module Queue(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [4:0] io_enq_bits_data,
  input  [1:0] io_enq_bits_dataType,
  input  [7:0] io_enq_bits_positon_col,
  input        io_deq_ready,
  output       io_deq_valid,
  output [4:0] io_deq_bits_data,
  output [1:0] io_deq_bits_dataType,
  output [7:0] io_deq_bits_positon_col
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] ram_data [0:15]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_data_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16]
  reg [1:0] ram_dataType [0:15]; // @[Decoupled.scala 218:16]
  wire [1:0] ram_dataType_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_dataType_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [1:0] ram_dataType_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_dataType_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_dataType_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_dataType_MPORT_en; // @[Decoupled.scala 218:16]
  reg [7:0] ram_positon_col [0:15]; // @[Decoupled.scala 218:16]
  wire [7:0] ram_positon_col_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_positon_col_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [7:0] ram_positon_col_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_positon_col_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_positon_col_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_positon_col_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] value; // @[Counter.scala 60:40]
  reg [3:0] value_1; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _value_T_1 = value + 4'h1; // @[Counter.scala 76:24]
  wire [3:0] _value_T_3 = value_1 + 4'h1; // @[Counter.scala 76:24]
  assign ram_data_io_deq_bits_MPORT_addr = value_1;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_dataType_io_deq_bits_MPORT_addr = value_1;
  assign ram_dataType_io_deq_bits_MPORT_data = ram_dataType[ram_dataType_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_dataType_MPORT_data = io_enq_bits_dataType;
  assign ram_dataType_MPORT_addr = value;
  assign ram_dataType_MPORT_mask = 1'h1;
  assign ram_dataType_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_positon_col_io_deq_bits_MPORT_addr = value_1;
  assign ram_positon_col_io_deq_bits_MPORT_data = ram_positon_col[ram_positon_col_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_positon_col_MPORT_data = io_enq_bits_positon_col;
  assign ram_positon_col_MPORT_addr = value;
  assign ram_positon_col_MPORT_mask = 1'h1;
  assign ram_positon_col_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_dataType = ram_dataType_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_positon_col = ram_positon_col_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_dataType_MPORT_en & ram_dataType_MPORT_mask) begin
      ram_dataType[ram_dataType_MPORT_addr] <= ram_dataType_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_positon_col_MPORT_en & ram_positon_col_MPORT_mask) begin
      ram_positon_col[ram_positon_col_MPORT_addr] <= ram_positon_col_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      value_1 <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_dataType[initvar] = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_positon_col[initvar] = _RAND_2[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Node(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_row,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType,
  output [7:0] io_dataPackageOut_bits_positon_col
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_row) == -8'sh1; // @[Node.scala 38:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_row) == 8'sh0; // @[Node.scala 40:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h0;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 39:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_positon_col = q_io_deq_bits_positon_col; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 41:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_1(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh1; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h1;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module SRAM(
  input         clock,
  input         io_we,
  input  [7:0]  io_addr,
  input  [63:0] io_din,
  output [63:0] io_dout,
  input         io_rstLowas
);
  wire  ram_clk; // @[ipSram.scala 29:19]
  wire  ram_rst_n; // @[ipSram.scala 29:19]
  wire  ram_cs_n; // @[ipSram.scala 29:19]
  wire  ram_wr_n; // @[ipSram.scala 29:19]
  wire [7:0] ram_rd_addr; // @[ipSram.scala 29:19]
  wire [7:0] ram_wr_addr; // @[ipSram.scala 29:19]
  wire [63:0] ram_data_in; // @[ipSram.scala 29:19]
  wire [63:0] ram_data_out; // @[ipSram.scala 29:19]
  DW_ram_r_w_s_dff ram ( // @[ipSram.scala 29:19]
    .clk(ram_clk),
    .rst_n(ram_rst_n),
    .cs_n(ram_cs_n),
    .wr_n(ram_wr_n),
    .rd_addr(ram_rd_addr),
    .wr_addr(ram_wr_addr),
    .data_in(ram_data_in),
    .data_out(ram_data_out)
  );
  assign io_dout = ram_data_out; // @[ipSram.scala 37:11]
  assign ram_clk = clock; // @[ipSram.scala 30:14]
  assign ram_rst_n = io_rstLowas; // @[ipSram.scala 31:16]
  assign ram_cs_n = 1'h0; // @[ipSram.scala 32:15]
  assign ram_wr_n = io_we; // @[ipSram.scala 33:15]
  assign ram_rd_addr = io_addr; // @[ipSram.scala 34:18]
  assign ram_wr_addr = io_addr; // @[ipSram.scala 35:18]
  assign ram_data_in = io_din; // @[ipSram.scala 36:18]
endmodule
module PECore(
  input         clock,
  input         reset,
  input  [1:0]  io_stateSW,
  input  [15:0] io_regConfig_ochannelNum,
  input  [15:0] io_regConfig_filterLen,
  output        io_filter_ready,
  input         io_filter_valid,
  input  [15:0] io_filter_bits,
  output        io_ifmap_ready,
  input         io_ifmap_valid,
  input  [15:0] io_ifmap_bits,
  output        io_pSumIn_ready,
  input         io_pSumIn_valid,
  input  [63:0] io_pSumIn_bits,
  input         io_pSumOut_ready,
  output        io_pSumOut_valid,
  output [63:0] io_pSumOut_bits,
  output [3:0]  io_stateOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  pSumSRAM_clock; // @[PECore.scala 48:26]
  wire  pSumSRAM_io_we; // @[PECore.scala 48:26]
  wire [7:0] pSumSRAM_io_addr; // @[PECore.scala 48:26]
  wire [63:0] pSumSRAM_io_din; // @[PECore.scala 48:26]
  wire [63:0] pSumSRAM_io_dout; // @[PECore.scala 48:26]
  wire  pSumSRAM_io_rstLowas; // @[PECore.scala 48:26]
  reg [1:0] state; // @[PECore.scala 53:24]
  reg [10:0] value; // @[Counter.scala 60:40]
  reg [7:0] value_1; // @[Counter.scala 60:40]
  reg [7:0] value_3; // @[Counter.scala 60:40]
  wire [15:0] _GEN_63 = {{8'd0}, value_1}; // @[PECore.scala 65:58]
  wire  clrDone = state == 2'h0 & _GEN_63 == io_regConfig_ochannelNum; // @[PECore.scala 65:43]
  wire [31:0] _T_6 = $signed(io_filter_bits) * $signed(io_ifmap_bits); // @[PECore.scala 78:40]
  wire [63:0] _GEN_64 = {{32{_T_6[31]}},_T_6}; // @[PECore.scala 78:56]
  wire [63:0] pRes = $signed(_GEN_64) + $signed(pSumSRAM_io_dout); // @[PECore.scala 78:56]
  wire  _T_11 = io_filter_ready & io_filter_valid; // @[Decoupled.scala 40:37]
  wire  _T_15 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire [7:0] _value_T_1 = value_1 + 8'h1; // @[Counter.scala 76:24]
  wire [7:0] _GEN_2 = _GEN_63 < io_regConfig_ochannelNum ? value_1 : value_3; // @[PECore.scala 104:55 ipSram.scala 45:13 ipSram.scala 40:13]
  wire  _GEN_3 = _GEN_63 < io_regConfig_ochannelNum ? 1'h0 : 1'h1; // @[PECore.scala 104:55 ipSram.scala 46:11 ipSram.scala 41:11]
  wire  _T_19 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [15:0] _T_24 = io_regConfig_filterLen - 16'h1; // @[PECore.scala 115:59]
  wire [15:0] _GEN_66 = {{5'd0}, value}; // @[PECore.scala 115:35]
  wire  _T_25 = _GEN_66 == _T_24; // @[PECore.scala 115:35]
  wire [1:0] _GEN_5 = _GEN_66 == _T_24 ? 2'h2 : state; // @[PECore.scala 115:66 PECore.scala 116:27 PECore.scala 53:24]
  wire [10:0] _value_T_3 = value + 11'h1; // @[Counter.scala 76:24]
  wire [10:0] _GEN_6 = _T_25 ? 11'h0 : _value_T_3; // @[PECore.scala 118:66 PECore.scala 119:34 Counter.scala 76:15]
  wire [15:0] _T_30 = io_regConfig_ochannelNum - 16'h1; // @[PECore.scala 124:66]
  wire [15:0] _GEN_68 = {{8'd0}, value_3}; // @[PECore.scala 124:40]
  wire  _T_31 = _GEN_68 == _T_30; // @[PECore.scala 124:40]
  wire [7:0] _value_T_7 = value_3 + 8'h1; // @[Counter.scala 76:24]
  wire [7:0] _GEN_8 = _GEN_68 == _T_30 ? 8'h0 : _value_T_7; // @[PECore.scala 124:72 PECore.scala 125:39 Counter.scala 76:15]
  wire  _GEN_12 = _T_11 & io_ifmap_valid ? 1'h0 : 1'h1; // @[PECore.scala 112:61 ipSram.scala 46:11 ipSram.scala 41:11]
  wire [63:0] _GEN_13 = _T_11 & io_ifmap_valid ? $signed(pRes) : $signed(64'sh0); // @[PECore.scala 112:61 ipSram.scala 47:12 PECore.scala 50:21]
  wire  _GEN_17 = _T_11 & io_ifmap_valid & _T_31; // @[PECore.scala 112:61 PECore.scala 70:20]
  wire  _T_35 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_36 = io_pSumIn_ready & io_pSumIn_valid; // @[Decoupled.scala 40:37]
  wire  _T_38 = _T_36 & io_pSumOut_ready; // @[PECore.scala 140:35]
  wire [1:0] _GEN_20 = _T_31 ? 2'h3 : state; // @[PECore.scala 142:72 PECore.scala 144:27 PECore.scala 53:24]
  wire [63:0] _T_44 = $signed(pSumSRAM_io_dout) + $signed(io_pSumIn_bits); // @[PECore.scala 148:65]
  wire [7:0] _GEN_21 = _T_36 & io_pSumOut_ready ? _GEN_8 : 8'h0; // @[PECore.scala 140:63 PECore.scala 138:31]
  wire [1:0] _GEN_22 = _T_36 & io_pSumOut_ready ? _GEN_20 : state; // @[PECore.scala 140:63 PECore.scala 53:24]
  wire [63:0] _GEN_25 = _T_36 & io_pSumOut_ready ? $signed(_T_44) : $signed(64'sh0); // @[PECore.scala 140:63 PECore.scala 148:33 PECore.scala 73:21]
  wire  _T_45 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_27 = _T_45 ? 8'h0 : value_1; // @[Conditional.scala 39:67 PECore.scala 154:26 Counter.scala 60:40]
  wire [1:0] _GEN_28 = _T_45 ? 2'h0 : state; // @[Conditional.scala 39:67 PECore.scala 160:19 PECore.scala 53:24]
  wire [63:0] _GEN_34 = _T_35 ? $signed(_GEN_25) : $signed(64'sh0); // @[Conditional.scala 39:67 PECore.scala 73:21]
  wire  _GEN_39 = _T_19 ? _GEN_12 : 1'h1; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_40 = _T_19 ? $signed(_GEN_13) : $signed(64'sh0); // @[Conditional.scala 39:67 PECore.scala 50:21]
  wire  _GEN_44 = _T_19 & _GEN_17; // @[Conditional.scala 39:67 PECore.scala 70:20]
  wire  _GEN_46 = _T_19 ? 1'h0 : _T_35; // @[Conditional.scala 39:67 PECore.scala 68:21]
  wire [63:0] _GEN_47 = _T_19 ? $signed(64'sh0) : $signed(_GEN_34); // @[Conditional.scala 39:67 PECore.scala 73:21]
  wire  _GEN_48 = _T_19 ? 1'h0 : _T_35 & _T_38; // @[Conditional.scala 39:67 PECore.scala 72:22]
  SRAM pSumSRAM ( // @[PECore.scala 48:26]
    .clock(pSumSRAM_clock),
    .io_we(pSumSRAM_io_we),
    .io_addr(pSumSRAM_io_addr),
    .io_din(pSumSRAM_io_din),
    .io_dout(pSumSRAM_io_dout),
    .io_rstLowas(pSumSRAM_io_rstLowas)
  );
  assign io_filter_ready = _T_15 ? 1'h0 : _T_19; // @[Conditional.scala 40:58 PECore.scala 69:21]
  assign io_ifmap_ready = _T_15 ? 1'h0 : _GEN_44; // @[Conditional.scala 40:58 PECore.scala 70:20]
  assign io_pSumIn_ready = _T_15 ? 1'h0 : _GEN_46; // @[Conditional.scala 40:58 PECore.scala 68:21]
  assign io_pSumOut_valid = _T_15 ? 1'h0 : _GEN_48; // @[Conditional.scala 40:58 PECore.scala 72:22]
  assign io_pSumOut_bits = _T_15 ? $signed(64'sh0) : $signed(_GEN_47); // @[Conditional.scala 40:58 PECore.scala 73:21]
  assign io_stateOut = {{2'd0}, state}; // @[PECore.scala 75:17]
  assign pSumSRAM_clock = clock;
  assign pSumSRAM_io_we = _T_15 ? _GEN_3 : _GEN_39; // @[Conditional.scala 40:58]
  assign pSumSRAM_io_addr = _T_15 ? _GEN_2 : value_3; // @[Conditional.scala 40:58]
  assign pSumSRAM_io_din = _T_15 ? $signed(64'sh0) : $signed(_GEN_40); // @[Conditional.scala 40:58]
  assign pSumSRAM_io_rstLowas = reset + 1'h1; // @[PECore.scala 49:44]
  always @(posedge clock) begin
    if (reset) begin // @[PECore.scala 53:24]
      state <= 2'h0; // @[PECore.scala 53:24]
    end else if (_T_15) begin // @[Conditional.scala 40:58]
      if (io_stateSW == 2'h1 & clrDone) begin // @[PECore.scala 100:48]
        state <= 2'h1; // @[PECore.scala 101:23]
      end
    end else if (_T_19) begin // @[Conditional.scala 39:67]
      if (_T_11 & io_ifmap_valid) begin // @[PECore.scala 112:61]
        state <= _GEN_5;
      end
    end else if (_T_35) begin // @[Conditional.scala 39:67]
      state <= _GEN_22;
    end else begin
      state <= _GEN_28;
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 11'h0; // @[Counter.scala 60:40]
    end else if (_T_15) begin // @[Conditional.scala 40:58]
      value <= 11'h0; // @[PECore.scala 91:26]
    end else if (_T_19) begin // @[Conditional.scala 39:67]
      if (_T_11 & io_ifmap_valid) begin // @[PECore.scala 112:61]
        value <= _GEN_6;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 8'h0; // @[Counter.scala 60:40]
    end else if (_T_15) begin // @[Conditional.scala 40:58]
      if (_GEN_63 < io_regConfig_ochannelNum) begin // @[PECore.scala 104:55]
        value_1 <= _value_T_1; // @[Counter.scala 76:15]
      end
    end else if (!(_T_19)) begin // @[Conditional.scala 39:67]
      if (!(_T_35)) begin // @[Conditional.scala 39:67]
        value_1 <= _GEN_27;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_3 <= 8'h0; // @[Counter.scala 60:40]
    end else if (_T_15) begin // @[Conditional.scala 40:58]
      value_3 <= 8'h0; // @[PECore.scala 94:31]
    end else if (_T_19) begin // @[Conditional.scala 39:67]
      if (_T_11 & io_ifmap_valid) begin // @[PECore.scala 112:61]
        value_3 <= _GEN_8;
      end
    end else if (_T_35) begin // @[Conditional.scala 39:67]
      value_3 <= _GEN_21;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  value_3 = _RAND_3[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_2(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] ram [0:2047]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [10:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_MPORT_data; // @[Decoupled.scala 218:16]
  wire [10:0] ram_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_en; // @[Decoupled.scala 218:16]
  reg [10:0] value; // @[Counter.scala 60:40]
  reg [10:0] value_1; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [10:0] _value_T_1 = value + 11'h1; // @[Counter.scala 76:24]
  wire [10:0] _value_T_3 = value_1 + 11'h1; // @[Counter.scala 76:24]
  assign ram_io_deq_bits_MPORT_addr = value_1;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 11'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 11'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      value_1 <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    ram[initvar] = _RAND_0[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[10:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_3(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [15:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [15:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] ram [0:255]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [7:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_MPORT_data; // @[Decoupled.scala 218:16]
  wire [7:0] ram_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_en; // @[Decoupled.scala 218:16]
  reg [7:0] value; // @[Counter.scala 60:40]
  reg [7:0] value_1; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [7:0] _value_T_1 = value + 8'h1; // @[Counter.scala 76:24]
  wire [7:0] _value_T_3 = value_1 + 8'h1; // @[Counter.scala 76:24]
  assign ram_io_deq_bits_MPORT_addr = value_1;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 8'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 8'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      value_1 <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_4(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram [0:255]; // @[Decoupled.scala 218:16]
  wire [63:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [7:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram_MPORT_data; // @[Decoupled.scala 218:16]
  wire [7:0] ram_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_en; // @[Decoupled.scala 218:16]
  reg [7:0] value; // @[Counter.scala 60:40]
  reg [7:0] value_1; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [7:0] _value_T_1 = value + 8'h1; // @[Counter.scala 76:24]
  wire [7:0] _value_T_3 = value_1 + 8'h1; // @[Counter.scala 76:24]
  assign ram_io_deq_bits_MPORT_addr = value_1;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 8'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 8'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      value_1 <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE(
  input         clock,
  input         reset,
  input  [1:0]  io_stateSW,
  output        io_peconfig_ready,
  input         io_peconfig_valid,
  input  [15:0] io_peconfig_bits_ichannelNum,
  input  [15:0] io_peconfig_bits_ochannelNum,
  input  [15:0] io_peconfig_bits_ofmapW,
  input  [15:0] io_peconfig_bits_stepW,
  input  [15:0] io_peconfig_bits_filterLen,
  input  [15:0] io_peconfig_bits_ifmapLen,
  output        io_filter_ready,
  input         io_filter_valid,
  input  [15:0] io_filter_bits,
  output        io_ifmap_ready,
  input         io_ifmap_valid,
  input  [15:0] io_ifmap_bits,
  output        io_pSumIn_ready,
  input         io_pSumIn_valid,
  input  [63:0] io_pSumIn_bits,
  input         io_pSumOut_ready,
  output        io_pSumOut_valid,
  output [63:0] io_pSumOut_bits,
  output [3:0]  io_stateOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  pecore_clock; // @[PE.scala 26:22]
  wire  pecore_reset; // @[PE.scala 26:22]
  wire [1:0] pecore_io_stateSW; // @[PE.scala 26:22]
  wire [15:0] pecore_io_regConfig_ochannelNum; // @[PE.scala 26:22]
  wire [15:0] pecore_io_regConfig_filterLen; // @[PE.scala 26:22]
  wire  pecore_io_filter_ready; // @[PE.scala 26:22]
  wire  pecore_io_filter_valid; // @[PE.scala 26:22]
  wire [15:0] pecore_io_filter_bits; // @[PE.scala 26:22]
  wire  pecore_io_ifmap_ready; // @[PE.scala 26:22]
  wire  pecore_io_ifmap_valid; // @[PE.scala 26:22]
  wire [15:0] pecore_io_ifmap_bits; // @[PE.scala 26:22]
  wire  pecore_io_pSumIn_ready; // @[PE.scala 26:22]
  wire  pecore_io_pSumIn_valid; // @[PE.scala 26:22]
  wire [63:0] pecore_io_pSumIn_bits; // @[PE.scala 26:22]
  wire  pecore_io_pSumOut_ready; // @[PE.scala 26:22]
  wire  pecore_io_pSumOut_valid; // @[PE.scala 26:22]
  wire [63:0] pecore_io_pSumOut_bits; // @[PE.scala 26:22]
  wire [3:0] pecore_io_stateOut; // @[PE.scala 26:22]
  wire  fQIn_clock; // @[Decoupled.scala 296:21]
  wire  fQIn_reset; // @[Decoupled.scala 296:21]
  wire  fQIn_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  fQIn_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [15:0] fQIn_io_enq_bits; // @[Decoupled.scala 296:21]
  wire  fQIn_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  fQIn_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [15:0] fQIn_io_deq_bits; // @[Decoupled.scala 296:21]
  wire  iQIn_clock; // @[Decoupled.scala 296:21]
  wire  iQIn_reset; // @[Decoupled.scala 296:21]
  wire  iQIn_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  iQIn_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [15:0] iQIn_io_enq_bits; // @[Decoupled.scala 296:21]
  wire  iQIn_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  iQIn_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [15:0] iQIn_io_deq_bits; // @[Decoupled.scala 296:21]
  wire  pSumQIn_clock; // @[Decoupled.scala 296:21]
  wire  pSumQIn_reset; // @[Decoupled.scala 296:21]
  wire  pSumQIn_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  pSumQIn_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [63:0] pSumQIn_io_enq_bits; // @[Decoupled.scala 296:21]
  wire  pSumQIn_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  pSumQIn_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [63:0] pSumQIn_io_deq_bits; // @[Decoupled.scala 296:21]
  wire  oSumQOut_clock; // @[Decoupled.scala 296:21]
  wire  oSumQOut_reset; // @[Decoupled.scala 296:21]
  wire  oSumQOut_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  oSumQOut_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [63:0] oSumQOut_io_enq_bits; // @[Decoupled.scala 296:21]
  wire  oSumQOut_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  oSumQOut_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [63:0] oSumQOut_io_deq_bits; // @[Decoupled.scala 296:21]
  reg [2:0] state; // @[PE.scala 37:22]
  reg [15:0] configReg_ichannelNum; // @[PE.scala 40:22]
  reg [15:0] configReg_ochannelNum; // @[PE.scala 40:22]
  reg [15:0] configReg_ofmapW; // @[PE.scala 40:22]
  reg [15:0] configReg_stepW; // @[PE.scala 40:22]
  reg [15:0] configReg_filterLen; // @[PE.scala 40:22]
  reg [15:0] configReg_ifmapLen; // @[PE.scala 40:22]
  reg [2:0] pstateSWReg; // @[PE.scala 41:28]
  reg [7:0] value; // @[Counter.scala 60:40]
  reg [7:0] value_1; // @[Counter.scala 60:40]
  reg [10:0] value_2; // @[Counter.scala 60:40]
  wire [3:0] pstate = pecore_io_stateOut;
  wire  _T = pstate == 4'h1; // @[PE.scala 69:15]
  wire  _T_3 = pecore_io_ifmap_ready & pecore_io_ifmap_valid; // @[Decoupled.scala 40:37]
  wire  _T_5 = state == 3'h4; // @[PE.scala 79:37]
  wire  iQMuxIn_ready = iQIn_io_enq_ready; // @[PE.scala 23:21 Decoupled.scala 299:17]
  wire  _GEN_0 = (state == 3'h5 | state == 3'h4) & iQMuxIn_ready; // @[PE.scala 79:48 PE.scala 80:22 PE.scala 82:22]
  wire  _T_8 = pecore_io_filter_ready & pecore_io_filter_valid; // @[Decoupled.scala 40:37]
  wire  fQMuxIn_ready = fQIn_io_enq_ready; // @[PE.scala 24:21 Decoupled.scala 299:17]
  wire  _T_10 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_11 = io_peconfig_ready & io_peconfig_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_13 = io_ifmap_ready & io_ifmap_valid; // @[Decoupled.scala 40:37]
  wire [15:0] _T_15 = configReg_ifmapLen - 16'h1; // @[PE.scala 122:53]
  wire [15:0] _GEN_81 = {{5'd0}, value_2}; // @[PE.scala 122:31]
  wire [10:0] _value_T_1 = value_2 + 11'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_24 = _GEN_81 >= _T_15 ? 3'h1 : state; // @[PE.scala 122:60 PE.scala 123:17 PE.scala 37:22]
  wire [10:0] _GEN_25 = _GEN_81 >= _T_15 ? 11'h0 : _value_T_1; // @[PE.scala 122:60 PE.scala 124:28 Counter.scala 76:15]
  wire [2:0] _GEN_26 = _GEN_81 >= _T_15 ? 3'h1 : pstateSWReg; // @[PE.scala 122:60 PE.scala 125:23 PE.scala 41:28]
  wire  _T_17 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire [15:0] _T_20 = configReg_ofmapW - 16'h1; // @[PE.scala 137:47]
  wire [15:0] _GEN_82 = {{8'd0}, value}; // @[PE.scala 137:27]
  wire [7:0] _value_T_3 = value + 8'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_30 = _GEN_82 >= _T_20 ? 3'h6 : 3'h4; // @[PE.scala 137:54 PE.scala 138:17 PE.scala 140:17]
  wire [7:0] _GEN_31 = _GEN_82 >= _T_20 ? value : _value_T_3; // @[PE.scala 137:54 Counter.scala 60:40 Counter.scala 76:15]
  wire [7:0] _GEN_32 = pstate == 4'h3 ? 8'h0 : value_1; // @[PE.scala 134:30 PE.scala 135:24 Counter.scala 60:40]
  wire [2:0] _GEN_33 = pstate == 4'h3 ? 3'h0 : 3'h1; // @[PE.scala 134:30 PE.scala 136:21 PE.scala 133:19]
  wire [2:0] _GEN_34 = pstate == 4'h3 ? _GEN_30 : state; // @[PE.scala 134:30 PE.scala 37:22]
  wire [7:0] _GEN_35 = pstate == 4'h3 ? _GEN_31 : value; // @[PE.scala 134:30 Counter.scala 60:40]
  wire  _T_22 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_23 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_24 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [31:0] _T_26 = configReg_stepW * configReg_ichannelNum; // @[PE.scala 158:46]
  wire [31:0] _T_28 = _T_26 - 32'h1; // @[PE.scala 158:71]
  wire [31:0] _GEN_83 = {{24'd0}, value_1}; // @[PE.scala 158:26]
  wire  _T_29 = _GEN_83 >= _T_28; // @[PE.scala 158:26]
  wire [7:0] _value_T_5 = value_1 + 8'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_36 = _T_29 ? 3'h1 : state; // @[PE.scala 159:11 PE.scala 160:17 PE.scala 37:22]
  wire [7:0] _GEN_37 = _T_29 ? value_1 : _value_T_5; // @[PE.scala 159:11 Counter.scala 60:40 Counter.scala 76:15]
  wire [2:0] _GEN_38 = _T_13 ? _GEN_36 : state; // @[PE.scala 156:29 PE.scala 37:22]
  wire [7:0] _GEN_39 = _T_13 ? _GEN_37 : value_1; // @[PE.scala 156:29 Counter.scala 60:40]
  wire  _T_30 = 3'h6 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_84 = {{1'd0}, io_stateSW}; // @[PE.scala 168:23]
  wire [2:0] _GEN_40 = _GEN_84 == 3'h5 ? 3'h5 : state; // @[PE.scala 170:41 PE.scala 171:15 PE.scala 37:22]
  wire [2:0] _GEN_41 = _GEN_84 == 3'h0 ? 3'h0 : _GEN_40; // @[PE.scala 168:32 PE.scala 169:15]
  wire [2:0] _GEN_42 = _T_30 ? 3'h0 : pstateSWReg; // @[Conditional.scala 39:67 PE.scala 167:19 PE.scala 41:28]
  wire [2:0] _GEN_43 = _T_30 ? _GEN_41 : state; // @[Conditional.scala 39:67 PE.scala 37:22]
  wire [2:0] _GEN_44 = _T_24 ? 3'h0 : _GEN_42; // @[Conditional.scala 39:67 PE.scala 154:19]
  wire [2:0] _GEN_45 = _T_24 ? _GEN_38 : _GEN_43; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_46 = _T_24 ? _GEN_39 : value_1; // @[Conditional.scala 39:67 Counter.scala 60:40]
  wire [2:0] _GEN_47 = _T_23 ? 3'h0 : _GEN_45; // @[Conditional.scala 39:67 PE.scala 149:13]
  wire [2:0] _GEN_48 = _T_23 ? pstateSWReg : _GEN_44; // @[Conditional.scala 39:67 PE.scala 41:28]
  wire [7:0] _GEN_49 = _T_23 ? value_1 : _GEN_46; // @[Conditional.scala 39:67 Counter.scala 60:40]
  wire [2:0] _GEN_50 = _T_22 ? 3'h0 : _GEN_47; // @[Conditional.scala 39:67 PE.scala 146:13]
  wire [2:0] _GEN_51 = _T_22 ? pstateSWReg : _GEN_48; // @[Conditional.scala 39:67 PE.scala 41:28]
  wire [7:0] _GEN_52 = _T_22 ? value_1 : _GEN_49; // @[Conditional.scala 39:67 Counter.scala 60:40]
  PECore pecore ( // @[PE.scala 26:22]
    .clock(pecore_clock),
    .reset(pecore_reset),
    .io_stateSW(pecore_io_stateSW),
    .io_regConfig_ochannelNum(pecore_io_regConfig_ochannelNum),
    .io_regConfig_filterLen(pecore_io_regConfig_filterLen),
    .io_filter_ready(pecore_io_filter_ready),
    .io_filter_valid(pecore_io_filter_valid),
    .io_filter_bits(pecore_io_filter_bits),
    .io_ifmap_ready(pecore_io_ifmap_ready),
    .io_ifmap_valid(pecore_io_ifmap_valid),
    .io_ifmap_bits(pecore_io_ifmap_bits),
    .io_pSumIn_ready(pecore_io_pSumIn_ready),
    .io_pSumIn_valid(pecore_io_pSumIn_valid),
    .io_pSumIn_bits(pecore_io_pSumIn_bits),
    .io_pSumOut_ready(pecore_io_pSumOut_ready),
    .io_pSumOut_valid(pecore_io_pSumOut_valid),
    .io_pSumOut_bits(pecore_io_pSumOut_bits),
    .io_stateOut(pecore_io_stateOut)
  );
  Queue_2 fQIn ( // @[Decoupled.scala 296:21]
    .clock(fQIn_clock),
    .reset(fQIn_reset),
    .io_enq_ready(fQIn_io_enq_ready),
    .io_enq_valid(fQIn_io_enq_valid),
    .io_enq_bits(fQIn_io_enq_bits),
    .io_deq_ready(fQIn_io_deq_ready),
    .io_deq_valid(fQIn_io_deq_valid),
    .io_deq_bits(fQIn_io_deq_bits)
  );
  Queue_3 iQIn ( // @[Decoupled.scala 296:21]
    .clock(iQIn_clock),
    .reset(iQIn_reset),
    .io_enq_ready(iQIn_io_enq_ready),
    .io_enq_valid(iQIn_io_enq_valid),
    .io_enq_bits(iQIn_io_enq_bits),
    .io_deq_ready(iQIn_io_deq_ready),
    .io_deq_valid(iQIn_io_deq_valid),
    .io_deq_bits(iQIn_io_deq_bits)
  );
  Queue_4 pSumQIn ( // @[Decoupled.scala 296:21]
    .clock(pSumQIn_clock),
    .reset(pSumQIn_reset),
    .io_enq_ready(pSumQIn_io_enq_ready),
    .io_enq_valid(pSumQIn_io_enq_valid),
    .io_enq_bits(pSumQIn_io_enq_bits),
    .io_deq_ready(pSumQIn_io_deq_ready),
    .io_deq_valid(pSumQIn_io_deq_valid),
    .io_deq_bits(pSumQIn_io_deq_bits)
  );
  Queue_4 oSumQOut ( // @[Decoupled.scala 296:21]
    .clock(oSumQOut_clock),
    .reset(oSumQOut_reset),
    .io_enq_ready(oSumQOut_io_enq_ready),
    .io_enq_valid(oSumQOut_io_enq_valid),
    .io_enq_bits(oSumQOut_io_enq_bits),
    .io_deq_ready(oSumQOut_io_deq_ready),
    .io_deq_valid(oSumQOut_io_deq_valid),
    .io_deq_bits(oSumQOut_io_deq_bits)
  );
  assign io_peconfig_ready = 3'h0 == state; // @[Conditional.scala 37:30]
  assign io_filter_ready = _T ? 1'h0 : fQMuxIn_ready; // @[PE.scala 86:24 PE.scala 89:21 PE.scala 91:13]
  assign io_ifmap_ready = pstate == 4'h1 | state == 3'h1 ? 1'h0 : _GEN_0; // @[PE.scala 69:41 PE.scala 73:20]
  assign io_pSumIn_ready = pSumQIn_io_enq_ready; // @[Decoupled.scala 299:17]
  assign io_pSumOut_valid = oSumQOut_io_deq_valid; // @[PE.scala 58:12]
  assign io_pSumOut_bits = oSumQOut_io_deq_bits; // @[PE.scala 58:12]
  assign io_stateOut = {{1'd0}, state}; // @[PE.scala 66:15]
  assign pecore_clock = clock;
  assign pecore_reset = reset;
  assign pecore_io_stateSW = pstateSWReg[1:0]; // @[PE.scala 64:21]
  assign pecore_io_regConfig_ochannelNum = configReg_ochannelNum; // @[PE.scala 62:23]
  assign pecore_io_regConfig_filterLen = configReg_filterLen; // @[PE.scala 62:23]
  assign pecore_io_filter_valid = fQIn_io_deq_valid; // @[PE.scala 106:20]
  assign pecore_io_filter_bits = fQIn_io_deq_bits; // @[PE.scala 106:20]
  assign pecore_io_ifmap_valid = _T_5 ? 1'h0 : iQIn_io_deq_valid; // @[PE.scala 95:25 PE.scala 98:27 PE.scala 103:21]
  assign pecore_io_ifmap_bits = _T_5 ? $signed(16'sh0) : $signed(iQIn_io_deq_bits); // @[PE.scala 95:25 PE.scala 97:26 PE.scala 103:21]
  assign pecore_io_pSumIn_valid = pSumQIn_io_deq_valid; // @[PE.scala 63:20]
  assign pecore_io_pSumIn_bits = pSumQIn_io_deq_bits; // @[PE.scala 63:20]
  assign pecore_io_pSumOut_ready = oSumQOut_io_enq_ready; // @[Decoupled.scala 299:17]
  assign fQIn_clock = clock;
  assign fQIn_reset = reset;
  assign fQIn_io_enq_valid = _T ? _T_8 : io_filter_valid; // @[PE.scala 86:24 PE.scala 88:19 PE.scala 91:13]
  assign fQIn_io_enq_bits = _T ? $signed(pecore_io_filter_bits) : $signed(io_filter_bits); // @[PE.scala 86:24 PE.scala 87:18 PE.scala 91:13]
  assign fQIn_io_deq_ready = pecore_io_filter_ready; // @[PE.scala 106:20]
  assign iQIn_clock = clock;
  assign iQIn_reset = reset;
  assign iQIn_io_enq_valid = pstate == 4'h1 | state == 3'h1 ? _T_3 : io_ifmap_valid; // @[PE.scala 69:41 PE.scala 72:19 PE.scala 78:19]
  assign iQIn_io_enq_bits = pstate == 4'h1 | state == 3'h1 ? $signed(pecore_io_ifmap_bits) : $signed(io_ifmap_bits); // @[PE.scala 69:41 PE.scala 71:18 PE.scala 77:18]
  assign iQIn_io_deq_ready = _T_5 | pecore_io_ifmap_ready; // @[PE.scala 95:25 PE.scala 96:16 PE.scala 103:21]
  assign pSumQIn_clock = clock;
  assign pSumQIn_reset = reset;
  assign pSumQIn_io_enq_valid = io_pSumIn_valid; // @[Decoupled.scala 297:22]
  assign pSumQIn_io_enq_bits = io_pSumIn_bits; // @[Decoupled.scala 298:21]
  assign pSumQIn_io_deq_ready = pecore_io_pSumIn_ready; // @[PE.scala 63:20]
  assign oSumQOut_clock = clock;
  assign oSumQOut_reset = reset;
  assign oSumQOut_io_enq_valid = pecore_io_pSumOut_valid; // @[Decoupled.scala 297:22]
  assign oSumQOut_io_enq_bits = pecore_io_pSumOut_bits; // @[Decoupled.scala 298:21]
  assign oSumQOut_io_deq_ready = io_pSumOut_ready; // @[PE.scala 58:12]
  always @(posedge clock) begin
    if (reset) begin // @[PE.scala 37:22]
      state <= 3'h0; // @[PE.scala 37:22]
    end else if (_T_10) begin // @[Conditional.scala 40:58]
      if (_T_11) begin // @[PE.scala 111:32]
        state <= 3'h5; // @[PE.scala 113:15]
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (_T_13) begin // @[PE.scala 121:29]
        state <= _GEN_24;
      end
    end else if (_T_17) begin // @[Conditional.scala 39:67]
      state <= _GEN_34;
    end else begin
      state <= _GEN_50;
    end
    if (_T_10) begin // @[Conditional.scala 40:58]
      if (_T_11) begin // @[PE.scala 111:32]
        configReg_ichannelNum <= io_peconfig_bits_ichannelNum; // @[PE.scala 112:19]
      end
    end
    if (_T_10) begin // @[Conditional.scala 40:58]
      if (_T_11) begin // @[PE.scala 111:32]
        configReg_ochannelNum <= io_peconfig_bits_ochannelNum; // @[PE.scala 112:19]
      end
    end
    if (_T_10) begin // @[Conditional.scala 40:58]
      if (_T_11) begin // @[PE.scala 111:32]
        configReg_ofmapW <= io_peconfig_bits_ofmapW; // @[PE.scala 112:19]
      end
    end
    if (_T_10) begin // @[Conditional.scala 40:58]
      if (_T_11) begin // @[PE.scala 111:32]
        configReg_stepW <= io_peconfig_bits_stepW; // @[PE.scala 112:19]
      end
    end
    if (_T_10) begin // @[Conditional.scala 40:58]
      if (_T_11) begin // @[PE.scala 111:32]
        configReg_filterLen <= io_peconfig_bits_filterLen; // @[PE.scala 112:19]
      end
    end
    if (_T_10) begin // @[Conditional.scala 40:58]
      if (_T_11) begin // @[PE.scala 111:32]
        configReg_ifmapLen <= io_peconfig_bits_ifmapLen; // @[PE.scala 112:19]
      end
    end
    if (reset) begin // @[PE.scala 41:28]
      pstateSWReg <= 3'h0; // @[PE.scala 41:28]
    end else if (!(_T_10)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[PE.scala 121:29]
          pstateSWReg <= _GEN_26;
        end
      end else if (_T_17) begin // @[Conditional.scala 39:67]
        pstateSWReg <= _GEN_33;
      end else begin
        pstateSWReg <= _GEN_51;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 8'h0; // @[Counter.scala 60:40]
    end else if (!(_T_10)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          value <= _GEN_35;
        end
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 8'h0; // @[Counter.scala 60:40]
    end else if (!(_T_10)) begin // @[Conditional.scala 40:58]
      if (!(_T_12)) begin // @[Conditional.scala 39:67]
        if (_T_17) begin // @[Conditional.scala 39:67]
          value_1 <= _GEN_32;
        end else begin
          value_1 <= _GEN_52;
        end
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_2 <= 11'h0; // @[Counter.scala 60:40]
    end else if (!(_T_10)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (_T_13) begin // @[PE.scala 121:29]
          value_2 <= _GEN_25;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  configReg_ichannelNum = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  configReg_ochannelNum = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  configReg_ofmapW = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  configReg_stepW = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  configReg_filterLen = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  configReg_ifmapLen = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  pstateSWReg = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  value = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  value_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  value_2 = _RAND_10[10:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_6(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [4:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [4:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] ram [0:2047]; // @[Decoupled.scala 218:16]
  wire [4:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [10:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [4:0] ram_MPORT_data; // @[Decoupled.scala 218:16]
  wire [10:0] ram_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_en; // @[Decoupled.scala 218:16]
  reg [10:0] value; // @[Counter.scala 60:40]
  reg [10:0] value_1; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [10:0] _value_T_1 = value + 11'h1; // @[Counter.scala 76:24]
  wire [10:0] _value_T_3 = value_1 + 11'h1; // @[Counter.scala 76:24]
  assign ram_io_deq_bits_MPORT_addr = value_1;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 11'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 11'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      value_1 <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    ram[initvar] = _RAND_0[4:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[10:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_8(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [19:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [19:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [19:0] ram [0:2047]; // @[Decoupled.scala 218:16]
  wire [19:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [10:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [19:0] ram_MPORT_data; // @[Decoupled.scala 218:16]
  wire [10:0] ram_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_en; // @[Decoupled.scala 218:16]
  reg [10:0] value; // @[Counter.scala 60:40]
  reg [10:0] value_1; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [10:0] _value_T_1 = value + 11'h1; // @[Counter.scala 76:24]
  wire [10:0] _value_T_3 = value_1 + 11'h1; // @[Counter.scala 76:24]
  assign ram_io_deq_bits_MPORT_addr = value_1;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 11'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 11'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      value_1 <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    ram[initvar] = _RAND_0[19:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[10:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_9(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram [0:2047]; // @[Decoupled.scala 218:16]
  wire [63:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [10:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram_MPORT_data; // @[Decoupled.scala 218:16]
  wire [10:0] ram_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_en; // @[Decoupled.scala 218:16]
  reg [10:0] value; // @[Counter.scala 60:40]
  reg [10:0] value_1; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [10:0] _value_T_1 = value + 11'h1; // @[Counter.scala 76:24]
  wire [10:0] _value_T_3 = value_1 + 11'h1; // @[Counter.scala 76:24]
  assign ram_io_deq_bits_MPORT_addr = value_1;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 11'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 11'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      value_1 <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[10:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PETop(
  input         clock,
  input         reset,
  input  [1:0]  io_stateSW,
  output        io_peconfig_ready,
  input         io_peconfig_valid,
  input  [15:0] io_peconfig_bits_ichannelNum,
  input  [15:0] io_peconfig_bits_ochannelNum,
  input  [15:0] io_peconfig_bits_ofmapW,
  input  [15:0] io_peconfig_bits_stepW,
  input  [15:0] io_peconfig_bits_filterLen,
  input  [15:0] io_peconfig_bits_ifmapLen,
  output        io_filter_ready,
  input         io_filter_valid,
  input  [4:0]  io_filter_bits,
  output        io_ifmap_ready,
  input         io_ifmap_valid,
  input  [4:0]  io_ifmap_bits,
  output        io_pSumIn_ready,
  input         io_pSumIn_valid,
  input  [19:0] io_pSumIn_bits,
  input         io_pSumOut_ready,
  output        io_pSumOut_valid,
  output [19:0] io_pSumOut_bits,
  output [3:0]  io_stateOut
);
  wire  pe_clock; // @[PETop.scala 16:20]
  wire  pe_reset; // @[PETop.scala 16:20]
  wire [1:0] pe_io_stateSW; // @[PETop.scala 16:20]
  wire  pe_io_peconfig_ready; // @[PETop.scala 16:20]
  wire  pe_io_peconfig_valid; // @[PETop.scala 16:20]
  wire [15:0] pe_io_peconfig_bits_ichannelNum; // @[PETop.scala 16:20]
  wire [15:0] pe_io_peconfig_bits_ochannelNum; // @[PETop.scala 16:20]
  wire [15:0] pe_io_peconfig_bits_ofmapW; // @[PETop.scala 16:20]
  wire [15:0] pe_io_peconfig_bits_stepW; // @[PETop.scala 16:20]
  wire [15:0] pe_io_peconfig_bits_filterLen; // @[PETop.scala 16:20]
  wire [15:0] pe_io_peconfig_bits_ifmapLen; // @[PETop.scala 16:20]
  wire  pe_io_filter_ready; // @[PETop.scala 16:20]
  wire  pe_io_filter_valid; // @[PETop.scala 16:20]
  wire [15:0] pe_io_filter_bits; // @[PETop.scala 16:20]
  wire  pe_io_ifmap_ready; // @[PETop.scala 16:20]
  wire  pe_io_ifmap_valid; // @[PETop.scala 16:20]
  wire [15:0] pe_io_ifmap_bits; // @[PETop.scala 16:20]
  wire  pe_io_pSumIn_ready; // @[PETop.scala 16:20]
  wire  pe_io_pSumIn_valid; // @[PETop.scala 16:20]
  wire [63:0] pe_io_pSumIn_bits; // @[PETop.scala 16:20]
  wire  pe_io_pSumOut_ready; // @[PETop.scala 16:20]
  wire  pe_io_pSumOut_valid; // @[PETop.scala 16:20]
  wire [63:0] pe_io_pSumOut_bits; // @[PETop.scala 16:20]
  wire [3:0] pe_io_stateOut; // @[PETop.scala 16:20]
  wire  fIn_clock; // @[Decoupled.scala 296:21]
  wire  fIn_reset; // @[Decoupled.scala 296:21]
  wire  fIn_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  fIn_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] fIn_io_enq_bits; // @[Decoupled.scala 296:21]
  wire  fIn_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  fIn_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] fIn_io_deq_bits; // @[Decoupled.scala 296:21]
  wire  iIn_clock; // @[Decoupled.scala 296:21]
  wire  iIn_reset; // @[Decoupled.scala 296:21]
  wire  iIn_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  iIn_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] iIn_io_enq_bits; // @[Decoupled.scala 296:21]
  wire  iIn_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  iIn_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] iIn_io_deq_bits; // @[Decoupled.scala 296:21]
  wire  pSumIn_clock; // @[Decoupled.scala 296:21]
  wire  pSumIn_reset; // @[Decoupled.scala 296:21]
  wire  pSumIn_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  pSumIn_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [19:0] pSumIn_io_enq_bits; // @[Decoupled.scala 296:21]
  wire  pSumIn_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  pSumIn_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [19:0] pSumIn_io_deq_bits; // @[Decoupled.scala 296:21]
  wire  oSumOut2_clock; // @[Decoupled.scala 296:21]
  wire  oSumOut2_reset; // @[Decoupled.scala 296:21]
  wire  oSumOut2_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  oSumOut2_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [63:0] oSumOut2_io_enq_bits; // @[Decoupled.scala 296:21]
  wire  oSumOut2_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  oSumOut2_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [63:0] oSumOut2_io_deq_bits; // @[Decoupled.scala 296:21]
  PE pe ( // @[PETop.scala 16:20]
    .clock(pe_clock),
    .reset(pe_reset),
    .io_stateSW(pe_io_stateSW),
    .io_peconfig_ready(pe_io_peconfig_ready),
    .io_peconfig_valid(pe_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pe_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pe_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pe_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pe_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pe_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pe_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pe_io_filter_ready),
    .io_filter_valid(pe_io_filter_valid),
    .io_filter_bits(pe_io_filter_bits),
    .io_ifmap_ready(pe_io_ifmap_ready),
    .io_ifmap_valid(pe_io_ifmap_valid),
    .io_ifmap_bits(pe_io_ifmap_bits),
    .io_pSumIn_ready(pe_io_pSumIn_ready),
    .io_pSumIn_valid(pe_io_pSumIn_valid),
    .io_pSumIn_bits(pe_io_pSumIn_bits),
    .io_pSumOut_ready(pe_io_pSumOut_ready),
    .io_pSumOut_valid(pe_io_pSumOut_valid),
    .io_pSumOut_bits(pe_io_pSumOut_bits),
    .io_stateOut(pe_io_stateOut)
  );
  Queue_6 fIn ( // @[Decoupled.scala 296:21]
    .clock(fIn_clock),
    .reset(fIn_reset),
    .io_enq_ready(fIn_io_enq_ready),
    .io_enq_valid(fIn_io_enq_valid),
    .io_enq_bits(fIn_io_enq_bits),
    .io_deq_ready(fIn_io_deq_ready),
    .io_deq_valid(fIn_io_deq_valid),
    .io_deq_bits(fIn_io_deq_bits)
  );
  Queue_6 iIn ( // @[Decoupled.scala 296:21]
    .clock(iIn_clock),
    .reset(iIn_reset),
    .io_enq_ready(iIn_io_enq_ready),
    .io_enq_valid(iIn_io_enq_valid),
    .io_enq_bits(iIn_io_enq_bits),
    .io_deq_ready(iIn_io_deq_ready),
    .io_deq_valid(iIn_io_deq_valid),
    .io_deq_bits(iIn_io_deq_bits)
  );
  Queue_8 pSumIn ( // @[Decoupled.scala 296:21]
    .clock(pSumIn_clock),
    .reset(pSumIn_reset),
    .io_enq_ready(pSumIn_io_enq_ready),
    .io_enq_valid(pSumIn_io_enq_valid),
    .io_enq_bits(pSumIn_io_enq_bits),
    .io_deq_ready(pSumIn_io_deq_ready),
    .io_deq_valid(pSumIn_io_deq_valid),
    .io_deq_bits(pSumIn_io_deq_bits)
  );
  Queue_9 oSumOut2 ( // @[Decoupled.scala 296:21]
    .clock(oSumOut2_clock),
    .reset(oSumOut2_reset),
    .io_enq_ready(oSumOut2_io_enq_ready),
    .io_enq_valid(oSumOut2_io_enq_valid),
    .io_enq_bits(oSumOut2_io_enq_bits),
    .io_deq_ready(oSumOut2_io_deq_ready),
    .io_deq_valid(oSumOut2_io_deq_valid),
    .io_deq_bits(oSumOut2_io_deq_bits)
  );
  assign io_peconfig_ready = pe_io_peconfig_ready; // @[PETop.scala 27:20]
  assign io_filter_ready = fIn_io_enq_ready; // @[Decoupled.scala 299:17]
  assign io_ifmap_ready = iIn_io_enq_ready; // @[Decoupled.scala 299:17]
  assign io_pSumIn_ready = pSumIn_io_enq_ready; // @[Decoupled.scala 299:17]
  assign io_pSumOut_valid = oSumOut2_io_deq_valid; // @[PETop.scala 24:14]
  assign io_pSumOut_bits = oSumOut2_io_deq_bits[19:0]; // @[PETop.scala 24:14]
  assign io_stateOut = pe_io_stateOut; // @[PETop.scala 31:17]
  assign pe_clock = clock;
  assign pe_reset = reset;
  assign pe_io_stateSW = io_stateSW; // @[PETop.scala 29:19]
  assign pe_io_peconfig_valid = io_peconfig_valid; // @[PETop.scala 27:20]
  assign pe_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PETop.scala 27:20]
  assign pe_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PETop.scala 27:20]
  assign pe_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PETop.scala 27:20]
  assign pe_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PETop.scala 27:20]
  assign pe_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PETop.scala 27:20]
  assign pe_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PETop.scala 27:20]
  assign pe_io_filter_valid = fIn_io_deq_valid; // @[PETop.scala 25:18]
  assign pe_io_filter_bits = {{11{fIn_io_deq_bits[4]}},fIn_io_deq_bits}; // @[PETop.scala 25:18]
  assign pe_io_ifmap_valid = iIn_io_deq_valid; // @[PETop.scala 26:17]
  assign pe_io_ifmap_bits = {{11{iIn_io_deq_bits[4]}},iIn_io_deq_bits}; // @[PETop.scala 26:17]
  assign pe_io_pSumIn_valid = pSumIn_io_deq_valid; // @[PETop.scala 28:18]
  assign pe_io_pSumIn_bits = {{44{pSumIn_io_deq_bits[19]}},pSumIn_io_deq_bits}; // @[PETop.scala 28:18]
  assign pe_io_pSumOut_ready = oSumOut2_io_enq_ready; // @[Decoupled.scala 299:17]
  assign fIn_clock = clock;
  assign fIn_reset = reset;
  assign fIn_io_enq_valid = io_filter_valid; // @[Decoupled.scala 297:22]
  assign fIn_io_enq_bits = io_filter_bits; // @[Decoupled.scala 298:21]
  assign fIn_io_deq_ready = pe_io_filter_ready; // @[PETop.scala 25:18]
  assign iIn_clock = clock;
  assign iIn_reset = reset;
  assign iIn_io_enq_valid = io_ifmap_valid; // @[Decoupled.scala 297:22]
  assign iIn_io_enq_bits = io_ifmap_bits; // @[Decoupled.scala 298:21]
  assign iIn_io_deq_ready = pe_io_ifmap_ready; // @[PETop.scala 26:17]
  assign pSumIn_clock = clock;
  assign pSumIn_reset = reset;
  assign pSumIn_io_enq_valid = io_pSumIn_valid; // @[Decoupled.scala 297:22]
  assign pSumIn_io_enq_bits = io_pSumIn_bits; // @[Decoupled.scala 298:21]
  assign pSumIn_io_deq_ready = pe_io_pSumIn_ready; // @[PETop.scala 28:18]
  assign oSumOut2_clock = clock;
  assign oSumOut2_reset = reset;
  assign oSumOut2_io_enq_valid = pe_io_pSumOut_valid; // @[Decoupled.scala 297:22]
  assign oSumOut2_io_enq_bits = pe_io_pSumOut_bits; // @[Decoupled.scala 298:21]
  assign oSumOut2_io_deq_ready = io_pSumOut_ready; // @[PETop.scala 24:14]
endmodule
module dataSwitch(
  output        io_dataIn_ready,
  input         io_dataIn_valid,
  input  [15:0] io_dataIn_bits_data,
  input  [1:0]  io_dataIn_bits_dataType,
  input         io_filter_ready,
  output        io_filter_valid,
  output [15:0] io_filter_bits,
  input         io_ifmap_ready,
  output        io_ifmap_valid,
  output [15:0] io_ifmap_bits,
  input         io_pSum_ready,
  output        io_pSum_valid,
  output [15:0] io_pSum_bits
);
  wire [15:0] _GEN_0 = io_dataIn_bits_dataType == 2'h1 ? $signed(io_dataIn_bits_data) : $signed(16'sh0); // @[dataSwitch.scala 26:47 dataSwitch.scala 27:19 dataSwitch.scala 17:17]
  wire  _GEN_1 = io_dataIn_bits_dataType == 2'h1 & io_dataIn_valid; // @[dataSwitch.scala 26:47 dataSwitch.scala 28:20 dataSwitch.scala 18:18]
  wire  _GEN_2 = io_dataIn_bits_dataType == 2'h1 ? io_ifmap_ready : io_pSum_ready; // @[dataSwitch.scala 26:47 dataSwitch.scala 29:21 dataSwitch.scala 33:21]
  wire [15:0] _GEN_3 = io_dataIn_bits_dataType == 2'h1 ? $signed(16'sh0) : $signed(io_dataIn_bits_data); // @[dataSwitch.scala 26:47 dataSwitch.scala 19:16 dataSwitch.scala 31:18]
  wire  _GEN_4 = io_dataIn_bits_dataType == 2'h1 ? 1'h0 : io_dataIn_valid; // @[dataSwitch.scala 26:47 dataSwitch.scala 20:17 dataSwitch.scala 32:19]
  assign io_dataIn_ready = io_dataIn_bits_dataType == 2'h0 ? io_filter_ready : _GEN_2; // @[dataSwitch.scala 22:41 dataSwitch.scala 25:21]
  assign io_filter_valid = io_dataIn_bits_dataType == 2'h0 & io_dataIn_valid; // @[dataSwitch.scala 22:41 dataSwitch.scala 24:21 dataSwitch.scala 16:19]
  assign io_filter_bits = io_dataIn_bits_dataType == 2'h0 ? $signed(io_dataIn_bits_data) : $signed(16'sh0); // @[dataSwitch.scala 22:41 dataSwitch.scala 23:20 dataSwitch.scala 15:18]
  assign io_ifmap_valid = io_dataIn_bits_dataType == 2'h0 ? 1'h0 : _GEN_1; // @[dataSwitch.scala 22:41 dataSwitch.scala 18:18]
  assign io_ifmap_bits = io_dataIn_bits_dataType == 2'h0 ? $signed(16'sh0) : $signed(_GEN_0); // @[dataSwitch.scala 22:41 dataSwitch.scala 17:17]
  assign io_pSum_valid = io_dataIn_bits_dataType == 2'h0 ? 1'h0 : _GEN_4; // @[dataSwitch.scala 22:41 dataSwitch.scala 20:17]
  assign io_pSum_bits = io_dataIn_bits_dataType == 2'h0 ? $signed(16'sh0) : $signed(_GEN_3); // @[dataSwitch.scala 22:41 dataSwitch.scala 19:16]
endmodule
module Node_2(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh2; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h2;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_3(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh3; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h3;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_4(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh4; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h4;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_5(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh5; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h5;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_6(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh6; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h6;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_7(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh7; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h7;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_8(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh8; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h8;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_9(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh9; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h9;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_10(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sha; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'ha;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_11(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'shb; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'hb;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_12(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'shc; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'hc;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_13(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'shd; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'hd;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_14(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'she; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'he;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_15(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'shf; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'hf;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_16(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh10; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h10;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_17(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh11; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h11;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_18(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh12; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h12;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_19(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh13; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h13;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_20(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh14; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h14;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_21(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh15; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h15;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_22(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh16; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h16;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_23(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh17; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h17;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_24(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh18; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h0;
  wire [7:0] y = 8'h18;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_25(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_row,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType,
  output [7:0] io_dataPackageOut_bits_positon_col
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_row) == -8'sh1; // @[Node.scala 38:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_row) == 8'sh1; // @[Node.scala 40:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h0;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 39:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_positon_col = q_io_deq_bits_positon_col; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 41:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_26(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh1; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h1;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_27(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh2; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h2;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_28(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh3; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h3;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_29(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh4; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h4;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_30(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh5; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h5;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_31(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh6; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h6;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_32(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh7; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h7;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_33(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh8; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h8;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_34(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh9; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h9;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_35(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sha; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'ha;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_36(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'shb; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'hb;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_37(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'shc; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'hc;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_38(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'shd; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'hd;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_39(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'she; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'he;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_40(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'shf; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'hf;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_41(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh10; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h10;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_42(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh11; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h11;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_43(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh12; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h12;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_44(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh13; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h13;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_45(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh14; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h14;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_46(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh15; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h15;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_47(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh16; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h16;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_48(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh17; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h17;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_49(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh18; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h1;
  wire [7:0] y = 8'h18;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_50(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_row,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType,
  output [7:0] io_dataPackageOut_bits_positon_col
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_row) == -8'sh1; // @[Node.scala 38:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_row) == 8'sh2; // @[Node.scala 40:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h0;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 39:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_positon_col = q_io_deq_bits_positon_col; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 41:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_51(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh1; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h1;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_52(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh2; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h2;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_53(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh3; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h3;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_54(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh4; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h4;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_55(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh5; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h5;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_56(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh6; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h6;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_57(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh7; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h7;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_58(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh8; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h8;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_59(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh9; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h9;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_60(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sha; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'ha;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_61(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'shb; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'hb;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_62(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'shc; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'hc;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_63(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'shd; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'hd;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_64(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'she; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'he;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_65(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'shf; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'hf;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_66(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh10; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h10;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_67(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh11; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h11;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_68(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh12; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h12;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_69(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh13; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h13;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_70(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh14; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h14;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_71(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh15; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h15;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_72(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh16; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h16;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_73(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh17; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h17;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module Node_74(
  input        clock,
  input        reset,
  output       io_dataPackageIn_ready,
  input        io_dataPackageIn_valid,
  input  [4:0] io_dataPackageIn_bits_data,
  input  [1:0] io_dataPackageIn_bits_dataType,
  input  [7:0] io_dataPackageIn_bits_positon_col,
  input        io_dataPackageOut_ready,
  output       io_dataPackageOut_valid,
  output [4:0] io_dataPackageOut_bits_data,
  output [1:0] io_dataPackageOut_bits_dataType
);
  wire  q_clock; // @[Decoupled.scala 296:21]
  wire  q_reset; // @[Decoupled.scala 296:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_enq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_enq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_enq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 296:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 296:21]
  wire [4:0] q_io_deq_bits_data; // @[Decoupled.scala 296:21]
  wire [1:0] q_io_deq_bits_dataType; // @[Decoupled.scala 296:21]
  wire [7:0] q_io_deq_bits_positon_col; // @[Decoupled.scala 296:21]
  wire  boardcast = $signed(io_dataPackageIn_bits_positon_col) == -8'sh1; // @[Node.scala 44:53]
  wire  _T_2 = boardcast | $signed(io_dataPackageIn_bits_positon_col) == 8'sh18; // @[Node.scala 46:18]
  wire  qIn_ready = q_io_enq_ready; // @[Node.scala 29:17 Decoupled.scala 299:17]
  wire [7:0] x = 8'h2;
  wire [7:0] y = 8'h18;
  Queue q ( // @[Decoupled.scala 296:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_dataType(q_io_enq_bits_dataType),
    .io_enq_bits_positon_col(q_io_enq_bits_positon_col),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_dataType(q_io_deq_bits_dataType),
    .io_deq_bits_positon_col(q_io_deq_bits_positon_col)
  );
  assign io_dataPackageIn_ready = qIn_ready & _T_2; // @[Node.scala 45:41]
  assign io_dataPackageOut_valid = q_io_deq_valid; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_data = q_io_deq_bits_data; // @[Node.scala 33:5]
  assign io_dataPackageOut_bits_dataType = q_io_deq_bits_dataType; // @[Node.scala 33:5]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_dataPackageIn_valid & _T_2; // @[Node.scala 47:41]
  assign q_io_enq_bits_data = io_dataPackageIn_bits_data; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_dataType = io_dataPackageIn_bits_dataType; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_enq_bits_positon_col = io_dataPackageIn_bits_positon_col; // @[Node.scala 29:17 Node.scala 32:7]
  assign q_io_deq_ready = io_dataPackageOut_ready; // @[Node.scala 33:5]
endmodule
module PEArray(
  input         clock,
  input         reset,
  output        io_dataIn_ready,
  input         io_dataIn_valid,
  input  [4:0]  io_dataIn_bits_data,
  input  [1:0]  io_dataIn_bits_dataType,
  input  [7:0]  io_dataIn_bits_positon_row,
  input  [7:0]  io_dataIn_bits_positon_col,
  input  [1:0]  io_stateSW,
  output        io_peconfig_ready,
  input         io_peconfig_valid,
  input  [15:0] io_peconfig_bits_ichannelNum,
  input  [15:0] io_peconfig_bits_ochannelNum,
  input  [15:0] io_peconfig_bits_ifmapW,
  input  [15:0] io_peconfig_bits_ifmapH,
  input  [15:0] io_peconfig_bits_filterK,
  input  [15:0] io_peconfig_bits_ofmapW,
  input  [15:0] io_peconfig_bits_ofmapH,
  input  [15:0] io_peconfig_bits_stepW,
  input  [15:0] io_peconfig_bits_stepH,
  input  [15:0] io_peconfig_bits_filterLen,
  input  [15:0] io_peconfig_bits_ifmapLen,
  input         io_peconfig_bits_relu,
  input  [15:0] io_peconfig_bits_ID,
  input         io_oSumOut_0_ready,
  output        io_oSumOut_0_valid,
  output [19:0] io_oSumOut_0_bits,
  input         io_oSumOut_1_ready,
  output        io_oSumOut_1_valid,
  output [19:0] io_oSumOut_1_bits,
  input         io_oSumOut_2_ready,
  output        io_oSumOut_2_valid,
  output [19:0] io_oSumOut_2_bits,
  input         io_oSumOut_3_ready,
  output        io_oSumOut_3_valid,
  output [19:0] io_oSumOut_3_bits,
  input         io_oSumOut_4_ready,
  output        io_oSumOut_4_valid,
  output [19:0] io_oSumOut_4_bits,
  input         io_oSumOut_5_ready,
  output        io_oSumOut_5_valid,
  output [19:0] io_oSumOut_5_bits,
  input         io_oSumOut_6_ready,
  output        io_oSumOut_6_valid,
  output [19:0] io_oSumOut_6_bits,
  input         io_oSumOut_7_ready,
  output        io_oSumOut_7_valid,
  output [19:0] io_oSumOut_7_bits,
  input         io_oSumOut_8_ready,
  output        io_oSumOut_8_valid,
  output [19:0] io_oSumOut_8_bits,
  input         io_oSumOut_9_ready,
  output        io_oSumOut_9_valid,
  output [19:0] io_oSumOut_9_bits,
  input         io_oSumOut_10_ready,
  output        io_oSumOut_10_valid,
  output [19:0] io_oSumOut_10_bits,
  input         io_oSumOut_11_ready,
  output        io_oSumOut_11_valid,
  output [19:0] io_oSumOut_11_bits,
  input         io_oSumOut_12_ready,
  output        io_oSumOut_12_valid,
  output [19:0] io_oSumOut_12_bits,
  input         io_oSumOut_13_ready,
  output        io_oSumOut_13_valid,
  output [19:0] io_oSumOut_13_bits,
  input         io_oSumOut_14_ready,
  output        io_oSumOut_14_valid,
  output [19:0] io_oSumOut_14_bits,
  input         io_oSumOut_15_ready,
  output        io_oSumOut_15_valid,
  output [19:0] io_oSumOut_15_bits,
  input         io_oSumOut_16_ready,
  output        io_oSumOut_16_valid,
  output [19:0] io_oSumOut_16_bits,
  input         io_oSumOut_17_ready,
  output        io_oSumOut_17_valid,
  output [19:0] io_oSumOut_17_bits,
  input         io_oSumOut_18_ready,
  output        io_oSumOut_18_valid,
  output [19:0] io_oSumOut_18_bits,
  input         io_oSumOut_19_ready,
  output        io_oSumOut_19_valid,
  output [19:0] io_oSumOut_19_bits,
  input         io_oSumOut_20_ready,
  output        io_oSumOut_20_valid,
  output [19:0] io_oSumOut_20_bits,
  input         io_oSumOut_21_ready,
  output        io_oSumOut_21_valid,
  output [19:0] io_oSumOut_21_bits,
  input         io_oSumOut_22_ready,
  output        io_oSumOut_22_valid,
  output [19:0] io_oSumOut_22_bits,
  input         io_oSumOut_23_ready,
  output        io_oSumOut_23_valid,
  output [19:0] io_oSumOut_23_bits,
  output        io_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  NoC_0_0_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_0_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_0_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_0_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_0_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_0_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_0_io_dataPackageIn_bits_positon_row; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_0_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_0_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_1_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_1_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_1_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_1_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_1_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_1_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_1_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_1_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_1_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_1_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_1_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_0_clock; // @[PEArray.scala 36:24]
  wire  pes_0_0_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_0_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_0_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_0_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_0_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_0_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_0_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_0_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_0_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_0_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_0_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_0_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_0_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_0_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_0_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_0_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_0_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_0_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_0_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_0_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_0_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_0_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_0_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_0_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_0_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_0_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_0_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_0_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_0_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_0_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_0_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_0_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_0_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_0_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_0_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_0_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_2_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_2_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_2_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_2_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_2_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_2_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_2_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_2_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_2_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_2_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_2_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_1_clock; // @[PEArray.scala 36:24]
  wire  pes_0_1_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_1_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_1_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_1_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_1_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_1_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_1_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_1_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_1_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_1_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_1_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_1_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_1_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_1_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_1_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_1_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_1_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_1_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_1_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_1_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_1_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_1_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_1_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_1_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_1_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_1_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_1_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_1_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_1_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_1_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_1_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_1_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_1_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_1_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_1_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_1_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_3_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_3_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_3_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_3_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_3_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_3_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_3_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_3_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_3_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_3_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_3_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_2_clock; // @[PEArray.scala 36:24]
  wire  pes_0_2_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_2_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_2_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_2_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_2_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_2_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_2_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_2_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_2_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_2_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_2_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_2_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_2_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_2_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_2_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_2_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_2_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_2_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_2_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_2_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_2_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_2_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_2_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_2_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_2_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_2_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_2_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_2_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_2_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_2_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_2_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_2_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_2_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_2_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_2_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_2_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_4_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_4_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_4_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_4_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_4_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_4_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_4_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_4_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_4_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_4_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_4_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_3_clock; // @[PEArray.scala 36:24]
  wire  pes_0_3_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_3_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_3_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_3_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_3_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_3_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_3_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_3_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_3_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_3_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_3_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_3_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_3_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_3_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_3_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_3_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_3_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_3_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_3_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_3_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_3_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_3_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_3_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_3_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_3_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_3_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_3_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_3_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_3_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_3_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_3_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_3_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_3_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_3_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_3_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_3_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_5_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_5_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_5_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_5_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_5_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_5_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_5_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_5_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_5_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_5_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_5_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_4_clock; // @[PEArray.scala 36:24]
  wire  pes_0_4_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_4_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_4_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_4_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_4_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_4_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_4_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_4_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_4_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_4_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_4_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_4_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_4_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_4_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_4_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_4_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_4_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_4_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_4_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_4_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_4_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_4_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_4_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_4_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_4_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_4_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_4_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_4_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_4_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_4_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_4_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_4_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_4_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_4_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_4_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_4_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_6_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_6_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_6_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_6_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_6_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_6_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_6_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_6_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_6_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_6_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_6_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_5_clock; // @[PEArray.scala 36:24]
  wire  pes_0_5_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_5_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_5_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_5_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_5_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_5_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_5_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_5_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_5_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_5_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_5_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_5_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_5_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_5_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_5_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_5_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_5_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_5_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_5_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_5_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_5_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_5_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_5_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_5_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_5_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_5_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_5_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_5_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_5_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_5_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_5_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_5_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_5_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_5_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_5_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_5_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_7_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_7_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_7_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_7_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_7_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_7_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_7_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_7_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_7_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_7_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_7_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_6_clock; // @[PEArray.scala 36:24]
  wire  pes_0_6_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_6_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_6_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_6_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_6_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_6_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_6_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_6_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_6_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_6_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_6_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_6_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_6_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_6_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_6_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_6_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_6_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_6_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_6_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_6_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_6_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_6_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_6_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_6_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_6_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_6_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_6_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_6_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_6_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_6_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_6_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_6_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_6_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_6_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_6_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_6_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_8_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_8_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_8_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_8_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_8_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_8_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_8_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_8_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_8_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_8_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_8_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_7_clock; // @[PEArray.scala 36:24]
  wire  pes_0_7_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_7_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_7_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_7_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_7_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_7_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_7_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_7_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_7_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_7_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_7_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_7_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_7_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_7_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_7_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_7_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_7_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_7_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_7_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_7_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_7_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_7_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_7_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_7_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_7_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_7_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_7_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_7_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_7_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_7_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_7_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_7_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_7_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_7_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_7_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_7_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_9_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_9_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_9_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_9_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_9_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_9_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_9_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_9_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_9_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_9_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_9_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_8_clock; // @[PEArray.scala 36:24]
  wire  pes_0_8_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_8_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_8_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_8_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_8_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_8_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_8_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_8_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_8_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_8_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_8_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_8_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_8_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_8_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_8_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_8_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_8_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_8_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_8_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_8_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_8_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_8_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_8_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_8_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_8_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_8_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_8_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_8_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_8_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_8_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_8_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_8_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_8_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_8_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_8_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_8_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_10_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_10_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_10_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_10_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_10_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_10_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_10_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_10_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_10_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_10_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_10_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_9_clock; // @[PEArray.scala 36:24]
  wire  pes_0_9_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_9_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_9_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_9_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_9_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_9_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_9_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_9_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_9_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_9_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_9_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_9_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_9_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_9_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_9_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_9_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_9_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_9_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_9_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_9_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_9_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_9_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_9_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_9_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_9_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_9_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_9_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_9_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_9_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_9_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_9_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_9_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_9_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_9_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_9_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_9_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_11_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_11_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_11_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_11_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_11_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_11_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_11_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_11_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_11_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_11_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_11_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_10_clock; // @[PEArray.scala 36:24]
  wire  pes_0_10_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_10_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_10_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_10_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_10_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_10_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_10_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_10_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_10_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_10_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_10_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_10_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_10_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_10_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_10_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_10_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_10_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_10_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_10_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_10_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_10_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_10_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_10_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_10_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_10_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_10_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_10_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_10_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_10_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_10_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_10_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_10_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_10_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_10_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_10_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_10_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_12_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_12_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_12_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_12_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_12_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_12_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_12_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_12_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_12_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_12_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_12_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_11_clock; // @[PEArray.scala 36:24]
  wire  pes_0_11_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_11_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_11_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_11_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_11_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_11_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_11_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_11_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_11_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_11_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_11_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_11_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_11_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_11_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_11_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_11_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_11_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_11_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_11_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_11_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_11_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_11_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_11_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_11_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_11_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_11_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_11_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_11_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_11_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_11_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_11_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_11_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_11_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_11_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_11_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_11_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_13_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_13_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_13_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_13_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_13_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_13_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_13_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_13_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_13_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_13_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_13_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_12_clock; // @[PEArray.scala 36:24]
  wire  pes_0_12_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_12_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_12_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_12_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_12_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_12_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_12_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_12_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_12_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_12_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_12_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_12_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_12_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_12_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_12_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_12_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_12_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_12_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_12_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_12_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_12_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_12_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_12_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_12_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_12_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_12_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_12_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_12_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_12_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_12_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_12_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_12_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_12_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_12_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_12_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_12_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_14_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_14_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_14_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_14_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_14_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_14_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_14_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_14_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_14_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_14_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_14_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_13_clock; // @[PEArray.scala 36:24]
  wire  pes_0_13_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_13_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_13_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_13_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_13_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_13_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_13_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_13_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_13_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_13_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_13_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_13_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_13_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_13_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_13_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_13_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_13_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_13_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_13_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_13_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_13_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_13_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_13_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_13_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_13_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_13_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_13_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_13_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_13_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_13_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_13_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_13_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_13_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_13_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_13_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_13_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_15_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_15_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_15_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_15_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_15_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_15_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_15_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_15_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_15_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_15_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_15_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_14_clock; // @[PEArray.scala 36:24]
  wire  pes_0_14_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_14_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_14_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_14_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_14_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_14_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_14_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_14_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_14_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_14_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_14_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_14_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_14_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_14_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_14_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_14_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_14_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_14_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_14_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_14_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_14_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_14_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_14_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_14_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_14_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_14_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_14_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_14_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_14_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_14_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_14_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_14_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_14_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_14_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_14_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_14_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_16_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_16_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_16_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_16_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_16_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_16_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_16_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_16_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_16_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_16_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_16_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_15_clock; // @[PEArray.scala 36:24]
  wire  pes_0_15_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_15_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_15_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_15_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_15_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_15_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_15_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_15_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_15_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_15_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_15_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_15_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_15_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_15_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_15_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_15_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_15_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_15_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_15_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_15_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_15_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_15_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_15_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_15_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_15_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_15_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_15_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_15_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_15_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_15_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_15_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_15_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_15_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_15_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_15_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_15_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_17_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_17_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_17_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_17_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_17_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_17_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_17_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_17_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_17_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_17_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_17_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_16_clock; // @[PEArray.scala 36:24]
  wire  pes_0_16_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_16_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_16_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_16_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_16_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_16_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_16_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_16_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_16_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_16_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_16_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_16_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_16_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_16_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_16_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_16_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_16_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_16_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_16_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_16_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_16_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_16_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_16_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_16_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_16_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_16_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_16_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_16_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_16_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_16_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_16_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_16_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_16_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_16_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_16_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_16_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_18_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_18_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_18_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_18_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_18_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_18_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_18_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_18_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_18_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_18_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_18_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_17_clock; // @[PEArray.scala 36:24]
  wire  pes_0_17_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_17_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_17_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_17_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_17_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_17_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_17_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_17_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_17_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_17_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_17_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_17_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_17_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_17_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_17_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_17_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_17_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_17_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_17_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_17_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_17_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_17_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_17_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_17_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_17_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_17_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_17_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_17_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_17_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_17_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_17_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_17_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_17_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_17_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_17_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_17_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_19_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_19_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_19_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_19_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_19_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_19_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_19_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_19_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_19_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_19_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_19_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_18_clock; // @[PEArray.scala 36:24]
  wire  pes_0_18_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_18_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_18_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_18_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_18_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_18_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_18_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_18_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_18_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_18_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_18_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_18_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_18_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_18_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_18_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_18_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_18_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_18_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_18_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_18_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_18_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_18_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_18_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_18_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_18_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_18_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_18_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_18_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_18_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_18_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_18_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_18_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_18_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_18_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_18_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_18_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_20_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_20_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_20_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_20_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_20_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_20_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_20_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_20_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_20_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_20_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_20_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_19_clock; // @[PEArray.scala 36:24]
  wire  pes_0_19_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_19_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_19_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_19_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_19_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_19_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_19_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_19_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_19_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_19_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_19_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_19_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_19_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_19_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_19_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_19_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_19_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_19_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_19_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_19_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_19_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_19_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_19_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_19_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_19_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_19_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_19_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_19_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_19_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_19_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_19_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_19_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_19_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_19_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_19_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_19_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_21_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_21_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_21_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_21_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_21_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_21_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_21_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_21_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_21_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_21_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_21_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_20_clock; // @[PEArray.scala 36:24]
  wire  pes_0_20_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_20_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_20_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_20_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_20_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_20_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_20_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_20_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_20_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_20_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_20_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_20_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_20_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_20_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_20_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_20_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_20_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_20_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_20_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_20_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_20_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_20_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_20_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_20_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_20_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_20_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_20_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_20_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_20_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_20_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_20_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_20_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_20_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_20_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_20_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_20_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_22_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_22_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_22_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_22_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_22_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_22_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_22_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_22_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_22_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_22_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_22_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_21_clock; // @[PEArray.scala 36:24]
  wire  pes_0_21_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_21_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_21_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_21_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_21_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_21_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_21_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_21_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_21_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_21_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_21_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_21_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_21_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_21_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_21_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_21_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_21_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_21_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_21_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_21_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_21_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_21_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_21_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_21_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_21_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_21_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_21_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_21_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_21_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_21_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_21_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_21_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_21_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_21_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_21_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_21_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_23_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_23_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_23_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_23_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_23_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_23_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_23_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_23_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_23_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_23_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_23_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_22_clock; // @[PEArray.scala 36:24]
  wire  pes_0_22_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_22_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_22_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_22_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_22_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_22_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_22_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_22_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_22_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_22_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_22_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_22_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_22_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_22_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_22_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_22_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_22_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_22_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_22_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_22_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_22_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_22_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_22_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_22_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_22_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_22_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_22_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_22_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_22_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_22_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_22_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_22_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_22_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_22_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_22_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_22_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_0_24_clock; // @[PEArray.scala 34:24]
  wire  NoC_0_24_reset; // @[PEArray.scala 34:24]
  wire  NoC_0_24_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_24_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_24_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_24_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_0_24_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_0_24_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_0_24_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_0_24_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_0_24_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_0_23_clock; // @[PEArray.scala 36:24]
  wire  pes_0_23_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_0_23_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_0_23_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_0_23_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_23_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_23_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_23_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_23_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_23_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_0_23_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_0_23_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_0_23_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_23_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_0_23_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_0_23_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_0_23_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_0_23_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_0_23_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_23_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_0_23_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_0_23_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_0_23_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_0_23_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_0_23_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_0_23_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_23_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_0_23_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_0_23_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_0_23_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_23_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_0_23_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_0_23_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_23_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_0_23_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_0_23_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_0_23_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_0_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_0_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_0_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_0_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_0_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_0_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_0_io_dataPackageIn_bits_positon_row; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_0_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_0_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_1_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_1_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_1_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_1_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_1_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_1_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_1_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_1_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_1_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_1_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_1_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_0_clock; // @[PEArray.scala 36:24]
  wire  pes_1_0_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_0_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_0_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_0_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_0_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_0_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_0_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_0_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_0_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_0_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_0_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_0_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_0_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_0_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_0_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_0_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_0_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_0_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_0_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_0_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_0_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_0_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_0_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_0_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_0_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_0_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_0_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_0_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_0_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_0_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_0_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_0_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_0_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_0_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_0_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_0_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_2_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_2_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_2_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_2_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_2_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_2_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_2_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_2_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_2_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_2_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_2_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_1_clock; // @[PEArray.scala 36:24]
  wire  pes_1_1_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_1_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_1_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_1_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_1_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_1_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_1_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_1_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_1_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_1_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_1_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_1_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_1_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_1_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_1_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_1_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_1_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_1_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_1_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_1_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_1_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_1_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_1_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_1_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_1_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_1_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_1_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_1_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_1_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_1_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_1_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_1_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_1_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_1_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_1_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_1_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_3_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_3_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_3_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_3_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_3_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_3_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_3_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_3_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_3_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_3_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_3_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_2_clock; // @[PEArray.scala 36:24]
  wire  pes_1_2_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_2_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_2_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_2_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_2_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_2_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_2_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_2_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_2_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_2_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_2_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_2_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_2_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_2_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_2_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_2_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_2_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_2_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_2_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_2_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_2_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_2_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_2_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_2_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_2_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_2_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_2_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_2_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_2_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_2_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_2_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_2_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_2_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_2_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_2_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_2_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_4_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_4_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_4_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_4_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_4_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_4_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_4_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_4_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_4_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_4_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_4_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_3_clock; // @[PEArray.scala 36:24]
  wire  pes_1_3_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_3_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_3_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_3_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_3_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_3_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_3_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_3_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_3_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_3_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_3_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_3_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_3_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_3_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_3_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_3_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_3_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_3_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_3_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_3_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_3_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_3_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_3_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_3_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_3_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_3_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_3_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_3_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_3_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_3_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_3_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_3_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_3_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_3_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_3_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_3_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_5_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_5_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_5_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_5_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_5_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_5_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_5_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_5_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_5_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_5_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_5_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_4_clock; // @[PEArray.scala 36:24]
  wire  pes_1_4_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_4_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_4_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_4_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_4_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_4_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_4_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_4_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_4_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_4_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_4_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_4_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_4_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_4_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_4_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_4_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_4_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_4_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_4_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_4_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_4_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_4_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_4_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_4_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_4_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_4_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_4_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_4_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_4_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_4_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_4_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_4_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_4_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_4_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_4_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_4_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_6_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_6_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_6_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_6_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_6_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_6_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_6_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_6_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_6_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_6_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_6_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_5_clock; // @[PEArray.scala 36:24]
  wire  pes_1_5_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_5_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_5_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_5_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_5_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_5_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_5_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_5_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_5_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_5_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_5_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_5_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_5_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_5_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_5_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_5_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_5_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_5_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_5_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_5_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_5_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_5_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_5_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_5_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_5_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_5_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_5_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_5_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_5_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_5_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_5_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_5_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_5_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_5_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_5_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_5_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_7_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_7_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_7_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_7_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_7_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_7_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_7_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_7_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_7_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_7_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_7_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_6_clock; // @[PEArray.scala 36:24]
  wire  pes_1_6_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_6_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_6_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_6_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_6_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_6_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_6_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_6_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_6_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_6_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_6_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_6_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_6_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_6_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_6_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_6_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_6_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_6_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_6_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_6_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_6_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_6_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_6_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_6_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_6_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_6_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_6_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_6_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_6_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_6_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_6_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_6_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_6_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_6_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_6_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_6_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_8_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_8_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_8_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_8_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_8_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_8_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_8_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_8_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_8_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_8_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_8_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_7_clock; // @[PEArray.scala 36:24]
  wire  pes_1_7_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_7_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_7_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_7_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_7_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_7_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_7_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_7_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_7_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_7_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_7_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_7_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_7_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_7_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_7_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_7_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_7_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_7_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_7_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_7_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_7_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_7_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_7_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_7_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_7_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_7_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_7_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_7_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_7_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_7_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_7_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_7_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_7_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_7_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_7_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_7_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_9_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_9_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_9_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_9_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_9_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_9_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_9_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_9_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_9_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_9_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_9_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_8_clock; // @[PEArray.scala 36:24]
  wire  pes_1_8_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_8_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_8_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_8_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_8_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_8_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_8_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_8_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_8_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_8_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_8_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_8_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_8_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_8_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_8_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_8_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_8_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_8_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_8_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_8_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_8_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_8_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_8_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_8_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_8_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_8_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_8_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_8_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_8_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_8_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_8_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_8_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_8_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_8_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_8_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_8_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_10_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_10_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_10_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_10_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_10_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_10_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_10_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_10_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_10_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_10_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_10_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_9_clock; // @[PEArray.scala 36:24]
  wire  pes_1_9_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_9_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_9_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_9_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_9_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_9_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_9_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_9_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_9_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_9_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_9_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_9_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_9_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_9_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_9_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_9_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_9_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_9_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_9_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_9_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_9_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_9_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_9_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_9_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_9_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_9_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_9_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_9_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_9_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_9_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_9_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_9_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_9_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_9_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_9_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_9_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_11_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_11_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_11_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_11_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_11_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_11_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_11_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_11_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_11_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_11_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_11_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_10_clock; // @[PEArray.scala 36:24]
  wire  pes_1_10_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_10_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_10_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_10_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_10_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_10_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_10_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_10_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_10_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_10_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_10_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_10_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_10_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_10_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_10_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_10_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_10_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_10_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_10_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_10_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_10_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_10_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_10_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_10_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_10_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_10_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_10_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_10_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_10_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_10_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_10_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_10_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_10_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_10_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_10_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_10_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_12_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_12_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_12_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_12_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_12_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_12_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_12_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_12_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_12_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_12_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_12_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_11_clock; // @[PEArray.scala 36:24]
  wire  pes_1_11_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_11_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_11_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_11_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_11_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_11_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_11_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_11_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_11_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_11_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_11_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_11_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_11_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_11_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_11_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_11_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_11_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_11_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_11_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_11_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_11_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_11_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_11_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_11_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_11_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_11_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_11_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_11_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_11_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_11_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_11_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_11_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_11_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_11_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_11_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_11_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_13_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_13_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_13_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_13_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_13_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_13_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_13_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_13_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_13_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_13_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_13_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_12_clock; // @[PEArray.scala 36:24]
  wire  pes_1_12_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_12_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_12_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_12_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_12_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_12_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_12_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_12_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_12_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_12_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_12_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_12_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_12_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_12_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_12_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_12_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_12_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_12_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_12_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_12_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_12_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_12_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_12_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_12_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_12_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_12_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_12_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_12_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_12_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_12_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_12_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_12_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_12_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_12_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_12_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_12_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_14_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_14_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_14_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_14_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_14_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_14_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_14_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_14_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_14_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_14_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_14_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_13_clock; // @[PEArray.scala 36:24]
  wire  pes_1_13_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_13_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_13_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_13_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_13_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_13_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_13_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_13_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_13_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_13_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_13_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_13_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_13_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_13_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_13_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_13_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_13_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_13_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_13_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_13_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_13_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_13_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_13_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_13_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_13_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_13_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_13_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_13_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_13_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_13_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_13_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_13_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_13_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_13_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_13_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_13_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_15_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_15_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_15_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_15_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_15_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_15_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_15_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_15_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_15_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_15_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_15_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_14_clock; // @[PEArray.scala 36:24]
  wire  pes_1_14_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_14_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_14_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_14_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_14_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_14_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_14_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_14_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_14_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_14_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_14_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_14_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_14_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_14_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_14_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_14_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_14_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_14_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_14_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_14_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_14_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_14_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_14_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_14_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_14_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_14_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_14_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_14_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_14_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_14_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_14_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_14_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_14_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_14_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_14_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_14_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_16_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_16_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_16_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_16_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_16_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_16_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_16_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_16_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_16_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_16_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_16_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_15_clock; // @[PEArray.scala 36:24]
  wire  pes_1_15_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_15_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_15_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_15_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_15_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_15_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_15_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_15_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_15_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_15_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_15_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_15_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_15_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_15_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_15_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_15_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_15_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_15_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_15_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_15_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_15_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_15_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_15_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_15_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_15_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_15_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_15_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_15_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_15_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_15_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_15_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_15_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_15_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_15_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_15_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_15_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_17_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_17_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_17_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_17_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_17_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_17_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_17_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_17_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_17_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_17_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_17_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_16_clock; // @[PEArray.scala 36:24]
  wire  pes_1_16_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_16_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_16_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_16_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_16_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_16_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_16_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_16_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_16_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_16_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_16_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_16_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_16_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_16_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_16_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_16_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_16_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_16_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_16_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_16_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_16_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_16_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_16_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_16_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_16_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_16_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_16_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_16_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_16_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_16_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_16_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_16_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_16_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_16_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_16_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_16_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_18_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_18_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_18_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_18_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_18_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_18_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_18_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_18_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_18_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_18_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_18_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_17_clock; // @[PEArray.scala 36:24]
  wire  pes_1_17_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_17_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_17_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_17_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_17_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_17_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_17_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_17_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_17_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_17_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_17_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_17_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_17_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_17_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_17_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_17_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_17_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_17_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_17_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_17_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_17_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_17_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_17_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_17_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_17_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_17_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_17_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_17_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_17_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_17_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_17_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_17_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_17_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_17_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_17_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_17_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_19_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_19_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_19_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_19_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_19_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_19_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_19_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_19_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_19_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_19_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_19_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_18_clock; // @[PEArray.scala 36:24]
  wire  pes_1_18_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_18_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_18_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_18_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_18_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_18_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_18_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_18_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_18_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_18_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_18_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_18_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_18_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_18_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_18_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_18_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_18_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_18_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_18_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_18_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_18_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_18_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_18_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_18_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_18_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_18_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_18_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_18_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_18_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_18_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_18_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_18_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_18_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_18_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_18_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_18_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_20_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_20_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_20_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_20_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_20_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_20_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_20_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_20_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_20_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_20_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_20_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_19_clock; // @[PEArray.scala 36:24]
  wire  pes_1_19_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_19_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_19_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_19_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_19_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_19_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_19_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_19_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_19_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_19_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_19_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_19_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_19_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_19_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_19_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_19_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_19_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_19_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_19_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_19_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_19_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_19_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_19_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_19_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_19_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_19_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_19_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_19_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_19_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_19_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_19_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_19_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_19_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_19_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_19_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_19_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_21_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_21_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_21_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_21_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_21_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_21_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_21_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_21_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_21_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_21_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_21_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_20_clock; // @[PEArray.scala 36:24]
  wire  pes_1_20_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_20_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_20_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_20_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_20_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_20_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_20_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_20_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_20_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_20_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_20_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_20_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_20_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_20_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_20_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_20_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_20_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_20_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_20_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_20_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_20_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_20_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_20_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_20_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_20_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_20_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_20_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_20_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_20_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_20_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_20_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_20_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_20_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_20_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_20_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_20_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_22_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_22_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_22_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_22_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_22_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_22_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_22_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_22_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_22_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_22_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_22_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_21_clock; // @[PEArray.scala 36:24]
  wire  pes_1_21_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_21_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_21_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_21_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_21_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_21_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_21_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_21_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_21_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_21_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_21_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_21_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_21_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_21_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_21_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_21_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_21_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_21_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_21_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_21_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_21_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_21_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_21_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_21_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_21_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_21_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_21_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_21_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_21_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_21_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_21_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_21_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_21_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_21_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_21_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_21_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_23_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_23_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_23_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_23_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_23_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_23_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_23_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_23_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_23_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_23_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_23_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_22_clock; // @[PEArray.scala 36:24]
  wire  pes_1_22_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_22_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_22_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_22_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_22_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_22_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_22_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_22_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_22_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_22_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_22_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_22_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_22_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_22_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_22_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_22_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_22_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_22_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_22_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_22_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_22_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_22_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_22_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_22_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_22_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_22_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_22_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_22_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_22_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_22_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_22_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_22_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_22_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_22_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_22_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_22_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_1_24_clock; // @[PEArray.scala 34:24]
  wire  NoC_1_24_reset; // @[PEArray.scala 34:24]
  wire  NoC_1_24_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_24_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_24_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_24_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_1_24_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_1_24_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_1_24_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_1_24_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_1_24_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_1_23_clock; // @[PEArray.scala 36:24]
  wire  pes_1_23_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_1_23_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_1_23_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_1_23_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_23_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_23_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_23_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_23_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_23_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_1_23_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_1_23_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_1_23_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_23_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_1_23_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_1_23_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_1_23_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_1_23_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_1_23_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_23_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_1_23_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_1_23_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_1_23_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_1_23_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_1_23_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_1_23_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_23_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_1_23_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_1_23_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_1_23_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_23_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_1_23_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_1_23_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_23_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_1_23_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_1_23_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_1_23_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_0_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_0_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_0_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_0_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_0_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_0_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_0_io_dataPackageIn_bits_positon_row; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_0_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_0_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_1_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_1_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_1_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_1_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_1_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_1_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_1_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_1_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_1_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_1_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_1_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_0_clock; // @[PEArray.scala 36:24]
  wire  pes_2_0_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_0_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_0_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_0_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_0_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_0_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_0_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_0_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_0_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_0_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_0_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_0_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_0_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_0_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_0_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_0_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_0_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_0_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_0_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_0_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_0_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_0_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_0_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_0_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_0_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_0_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_0_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_0_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_0_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_0_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_0_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_0_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_0_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_0_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_0_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_0_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_2_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_2_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_2_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_2_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_2_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_2_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_2_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_2_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_2_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_2_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_2_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_1_clock; // @[PEArray.scala 36:24]
  wire  pes_2_1_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_1_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_1_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_1_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_1_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_1_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_1_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_1_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_1_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_1_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_1_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_1_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_1_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_1_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_1_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_1_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_1_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_1_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_1_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_1_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_1_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_1_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_1_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_1_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_1_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_1_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_1_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_1_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_1_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_1_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_1_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_1_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_1_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_1_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_1_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_1_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_3_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_3_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_3_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_3_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_3_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_3_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_3_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_3_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_3_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_3_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_3_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_2_clock; // @[PEArray.scala 36:24]
  wire  pes_2_2_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_2_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_2_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_2_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_2_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_2_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_2_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_2_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_2_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_2_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_2_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_2_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_2_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_2_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_2_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_2_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_2_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_2_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_2_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_2_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_2_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_2_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_2_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_2_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_2_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_2_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_2_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_2_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_2_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_2_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_2_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_2_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_2_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_2_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_2_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_2_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_4_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_4_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_4_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_4_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_4_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_4_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_4_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_4_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_4_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_4_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_4_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_3_clock; // @[PEArray.scala 36:24]
  wire  pes_2_3_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_3_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_3_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_3_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_3_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_3_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_3_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_3_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_3_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_3_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_3_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_3_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_3_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_3_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_3_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_3_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_3_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_3_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_3_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_3_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_3_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_3_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_3_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_3_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_3_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_3_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_3_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_3_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_3_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_3_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_3_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_3_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_3_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_3_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_3_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_3_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_5_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_5_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_5_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_5_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_5_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_5_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_5_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_5_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_5_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_5_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_5_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_4_clock; // @[PEArray.scala 36:24]
  wire  pes_2_4_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_4_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_4_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_4_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_4_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_4_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_4_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_4_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_4_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_4_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_4_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_4_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_4_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_4_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_4_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_4_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_4_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_4_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_4_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_4_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_4_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_4_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_4_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_4_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_4_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_4_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_4_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_4_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_4_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_4_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_4_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_4_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_4_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_4_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_4_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_4_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_6_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_6_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_6_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_6_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_6_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_6_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_6_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_6_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_6_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_6_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_6_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_5_clock; // @[PEArray.scala 36:24]
  wire  pes_2_5_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_5_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_5_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_5_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_5_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_5_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_5_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_5_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_5_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_5_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_5_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_5_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_5_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_5_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_5_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_5_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_5_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_5_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_5_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_5_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_5_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_5_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_5_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_5_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_5_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_5_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_5_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_5_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_5_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_5_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_5_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_5_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_5_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_5_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_5_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_5_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_7_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_7_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_7_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_7_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_7_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_7_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_7_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_7_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_7_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_7_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_7_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_6_clock; // @[PEArray.scala 36:24]
  wire  pes_2_6_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_6_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_6_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_6_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_6_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_6_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_6_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_6_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_6_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_6_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_6_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_6_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_6_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_6_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_6_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_6_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_6_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_6_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_6_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_6_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_6_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_6_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_6_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_6_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_6_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_6_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_6_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_6_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_6_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_6_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_6_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_6_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_6_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_6_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_6_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_6_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_8_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_8_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_8_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_8_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_8_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_8_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_8_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_8_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_8_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_8_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_8_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_7_clock; // @[PEArray.scala 36:24]
  wire  pes_2_7_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_7_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_7_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_7_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_7_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_7_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_7_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_7_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_7_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_7_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_7_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_7_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_7_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_7_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_7_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_7_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_7_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_7_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_7_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_7_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_7_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_7_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_7_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_7_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_7_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_7_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_7_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_7_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_7_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_7_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_7_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_7_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_7_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_7_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_7_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_7_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_9_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_9_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_9_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_9_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_9_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_9_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_9_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_9_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_9_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_9_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_9_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_8_clock; // @[PEArray.scala 36:24]
  wire  pes_2_8_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_8_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_8_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_8_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_8_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_8_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_8_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_8_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_8_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_8_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_8_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_8_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_8_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_8_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_8_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_8_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_8_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_8_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_8_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_8_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_8_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_8_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_8_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_8_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_8_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_8_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_8_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_8_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_8_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_8_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_8_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_8_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_8_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_8_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_8_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_8_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_10_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_10_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_10_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_10_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_10_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_10_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_10_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_10_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_10_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_10_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_10_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_9_clock; // @[PEArray.scala 36:24]
  wire  pes_2_9_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_9_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_9_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_9_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_9_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_9_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_9_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_9_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_9_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_9_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_9_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_9_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_9_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_9_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_9_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_9_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_9_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_9_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_9_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_9_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_9_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_9_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_9_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_9_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_9_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_9_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_9_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_9_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_9_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_9_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_9_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_9_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_9_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_9_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_9_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_9_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_11_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_11_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_11_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_11_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_11_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_11_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_11_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_11_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_11_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_11_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_11_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_10_clock; // @[PEArray.scala 36:24]
  wire  pes_2_10_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_10_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_10_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_10_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_10_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_10_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_10_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_10_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_10_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_10_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_10_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_10_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_10_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_10_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_10_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_10_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_10_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_10_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_10_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_10_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_10_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_10_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_10_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_10_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_10_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_10_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_10_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_10_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_10_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_10_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_10_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_10_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_10_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_10_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_10_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_10_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_12_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_12_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_12_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_12_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_12_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_12_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_12_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_12_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_12_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_12_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_12_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_11_clock; // @[PEArray.scala 36:24]
  wire  pes_2_11_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_11_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_11_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_11_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_11_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_11_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_11_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_11_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_11_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_11_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_11_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_11_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_11_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_11_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_11_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_11_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_11_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_11_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_11_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_11_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_11_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_11_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_11_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_11_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_11_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_11_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_11_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_11_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_11_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_11_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_11_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_11_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_11_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_11_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_11_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_11_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_13_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_13_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_13_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_13_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_13_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_13_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_13_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_13_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_13_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_13_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_13_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_12_clock; // @[PEArray.scala 36:24]
  wire  pes_2_12_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_12_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_12_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_12_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_12_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_12_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_12_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_12_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_12_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_12_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_12_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_12_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_12_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_12_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_12_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_12_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_12_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_12_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_12_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_12_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_12_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_12_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_12_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_12_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_12_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_12_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_12_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_12_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_12_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_12_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_12_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_12_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_12_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_12_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_12_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_12_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_14_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_14_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_14_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_14_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_14_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_14_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_14_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_14_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_14_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_14_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_14_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_13_clock; // @[PEArray.scala 36:24]
  wire  pes_2_13_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_13_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_13_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_13_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_13_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_13_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_13_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_13_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_13_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_13_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_13_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_13_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_13_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_13_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_13_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_13_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_13_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_13_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_13_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_13_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_13_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_13_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_13_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_13_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_13_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_13_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_13_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_13_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_13_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_13_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_13_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_13_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_13_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_13_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_13_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_13_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_15_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_15_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_15_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_15_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_15_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_15_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_15_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_15_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_15_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_15_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_15_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_14_clock; // @[PEArray.scala 36:24]
  wire  pes_2_14_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_14_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_14_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_14_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_14_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_14_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_14_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_14_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_14_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_14_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_14_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_14_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_14_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_14_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_14_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_14_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_14_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_14_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_14_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_14_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_14_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_14_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_14_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_14_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_14_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_14_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_14_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_14_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_14_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_14_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_14_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_14_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_14_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_14_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_14_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_14_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_16_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_16_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_16_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_16_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_16_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_16_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_16_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_16_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_16_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_16_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_16_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_15_clock; // @[PEArray.scala 36:24]
  wire  pes_2_15_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_15_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_15_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_15_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_15_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_15_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_15_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_15_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_15_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_15_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_15_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_15_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_15_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_15_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_15_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_15_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_15_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_15_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_15_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_15_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_15_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_15_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_15_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_15_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_15_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_15_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_15_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_15_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_15_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_15_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_15_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_15_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_15_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_15_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_15_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_15_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_17_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_17_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_17_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_17_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_17_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_17_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_17_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_17_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_17_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_17_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_17_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_16_clock; // @[PEArray.scala 36:24]
  wire  pes_2_16_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_16_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_16_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_16_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_16_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_16_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_16_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_16_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_16_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_16_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_16_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_16_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_16_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_16_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_16_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_16_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_16_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_16_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_16_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_16_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_16_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_16_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_16_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_16_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_16_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_16_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_16_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_16_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_16_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_16_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_16_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_16_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_16_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_16_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_16_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_16_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_18_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_18_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_18_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_18_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_18_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_18_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_18_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_18_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_18_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_18_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_18_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_17_clock; // @[PEArray.scala 36:24]
  wire  pes_2_17_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_17_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_17_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_17_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_17_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_17_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_17_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_17_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_17_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_17_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_17_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_17_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_17_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_17_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_17_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_17_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_17_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_17_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_17_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_17_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_17_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_17_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_17_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_17_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_17_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_17_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_17_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_17_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_17_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_17_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_17_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_17_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_17_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_17_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_17_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_17_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_19_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_19_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_19_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_19_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_19_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_19_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_19_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_19_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_19_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_19_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_19_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_18_clock; // @[PEArray.scala 36:24]
  wire  pes_2_18_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_18_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_18_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_18_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_18_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_18_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_18_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_18_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_18_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_18_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_18_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_18_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_18_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_18_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_18_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_18_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_18_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_18_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_18_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_18_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_18_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_18_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_18_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_18_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_18_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_18_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_18_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_18_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_18_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_18_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_18_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_18_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_18_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_18_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_18_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_18_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_20_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_20_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_20_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_20_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_20_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_20_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_20_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_20_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_20_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_20_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_20_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_19_clock; // @[PEArray.scala 36:24]
  wire  pes_2_19_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_19_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_19_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_19_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_19_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_19_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_19_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_19_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_19_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_19_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_19_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_19_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_19_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_19_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_19_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_19_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_19_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_19_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_19_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_19_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_19_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_19_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_19_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_19_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_19_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_19_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_19_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_19_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_19_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_19_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_19_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_19_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_19_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_19_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_19_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_19_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_21_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_21_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_21_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_21_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_21_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_21_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_21_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_21_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_21_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_21_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_21_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_20_clock; // @[PEArray.scala 36:24]
  wire  pes_2_20_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_20_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_20_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_20_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_20_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_20_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_20_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_20_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_20_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_20_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_20_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_20_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_20_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_20_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_20_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_20_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_20_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_20_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_20_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_20_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_20_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_20_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_20_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_20_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_20_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_20_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_20_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_20_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_20_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_20_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_20_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_20_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_20_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_20_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_20_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_20_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_22_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_22_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_22_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_22_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_22_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_22_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_22_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_22_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_22_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_22_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_22_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_21_clock; // @[PEArray.scala 36:24]
  wire  pes_2_21_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_21_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_21_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_21_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_21_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_21_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_21_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_21_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_21_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_21_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_21_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_21_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_21_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_21_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_21_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_21_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_21_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_21_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_21_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_21_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_21_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_21_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_21_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_21_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_21_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_21_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_21_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_21_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_21_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_21_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_21_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_21_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_21_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_21_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_21_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_21_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_23_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_23_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_23_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_23_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_23_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_23_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_23_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_23_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_23_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_23_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_23_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_22_clock; // @[PEArray.scala 36:24]
  wire  pes_2_22_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_22_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_22_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_22_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_22_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_22_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_22_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_22_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_22_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_22_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_22_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_22_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_22_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_22_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_22_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_22_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_22_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_22_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_22_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_22_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_22_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_22_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_22_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_22_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_22_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_22_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_22_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_22_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_22_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_22_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_22_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_22_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_22_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_22_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_22_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_22_io_pSum_bits; // @[PEArray.scala 37:24]
  wire  NoC_2_24_clock; // @[PEArray.scala 34:24]
  wire  NoC_2_24_reset; // @[PEArray.scala 34:24]
  wire  NoC_2_24_io_dataPackageIn_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_24_io_dataPackageIn_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_24_io_dataPackageIn_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_24_io_dataPackageIn_bits_dataType; // @[PEArray.scala 34:24]
  wire [7:0] NoC_2_24_io_dataPackageIn_bits_positon_col; // @[PEArray.scala 34:24]
  wire  NoC_2_24_io_dataPackageOut_ready; // @[PEArray.scala 34:24]
  wire  NoC_2_24_io_dataPackageOut_valid; // @[PEArray.scala 34:24]
  wire [4:0] NoC_2_24_io_dataPackageOut_bits_data; // @[PEArray.scala 34:24]
  wire [1:0] NoC_2_24_io_dataPackageOut_bits_dataType; // @[PEArray.scala 34:24]
  wire  pes_2_23_clock; // @[PEArray.scala 36:24]
  wire  pes_2_23_reset; // @[PEArray.scala 36:24]
  wire [1:0] pes_2_23_io_stateSW; // @[PEArray.scala 36:24]
  wire  pes_2_23_io_peconfig_ready; // @[PEArray.scala 36:24]
  wire  pes_2_23_io_peconfig_valid; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_23_io_peconfig_bits_ichannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_23_io_peconfig_bits_ochannelNum; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_23_io_peconfig_bits_ofmapW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_23_io_peconfig_bits_stepW; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_23_io_peconfig_bits_filterLen; // @[PEArray.scala 36:24]
  wire [15:0] pes_2_23_io_peconfig_bits_ifmapLen; // @[PEArray.scala 36:24]
  wire  pes_2_23_io_filter_ready; // @[PEArray.scala 36:24]
  wire  pes_2_23_io_filter_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_23_io_filter_bits; // @[PEArray.scala 36:24]
  wire  pes_2_23_io_ifmap_ready; // @[PEArray.scala 36:24]
  wire  pes_2_23_io_ifmap_valid; // @[PEArray.scala 36:24]
  wire [4:0] pes_2_23_io_ifmap_bits; // @[PEArray.scala 36:24]
  wire  pes_2_23_io_pSumIn_ready; // @[PEArray.scala 36:24]
  wire  pes_2_23_io_pSumIn_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_23_io_pSumIn_bits; // @[PEArray.scala 36:24]
  wire  pes_2_23_io_pSumOut_ready; // @[PEArray.scala 36:24]
  wire  pes_2_23_io_pSumOut_valid; // @[PEArray.scala 36:24]
  wire [19:0] pes_2_23_io_pSumOut_bits; // @[PEArray.scala 36:24]
  wire [3:0] pes_2_23_io_stateOut; // @[PEArray.scala 36:24]
  wire  dss_2_23_io_dataIn_ready; // @[PEArray.scala 37:24]
  wire  dss_2_23_io_dataIn_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_23_io_dataIn_bits_data; // @[PEArray.scala 37:24]
  wire [1:0] dss_2_23_io_dataIn_bits_dataType; // @[PEArray.scala 37:24]
  wire  dss_2_23_io_filter_ready; // @[PEArray.scala 37:24]
  wire  dss_2_23_io_filter_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_23_io_filter_bits; // @[PEArray.scala 37:24]
  wire  dss_2_23_io_ifmap_ready; // @[PEArray.scala 37:24]
  wire  dss_2_23_io_ifmap_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_23_io_ifmap_bits; // @[PEArray.scala 37:24]
  wire  dss_2_23_io_pSum_ready; // @[PEArray.scala 37:24]
  wire  dss_2_23_io_pSum_valid; // @[PEArray.scala 37:24]
  wire [15:0] dss_2_23_io_pSum_bits; // @[PEArray.scala 37:24]
  reg  doneReg; // @[PEArray.scala 17:24]
  reg  configReg_relu; // @[PEArray.scala 20:22]
  wire  _T = io_peconfig_ready & io_peconfig_valid; // @[Decoupled.scala 40:37]
  wire  _T_159 = pes_2_15_io_stateOut == 4'h6; // @[PEArray.scala 103:48]
  wire  _T_182 = pes_2_0_io_stateOut == 4'h6 | pes_2_1_io_stateOut == 4'h6 | pes_2_2_io_stateOut == 4'h6 |
    pes_2_3_io_stateOut == 4'h6 | pes_2_4_io_stateOut == 4'h6 | pes_2_5_io_stateOut == 4'h6 | pes_2_6_io_stateOut == 4'h6
     | pes_2_7_io_stateOut == 4'h6 | pes_2_8_io_stateOut == 4'h6 | pes_2_9_io_stateOut == 4'h6 | pes_2_10_io_stateOut
     == 4'h6 | pes_2_11_io_stateOut == 4'h6 | pes_2_12_io_stateOut == 4'h6 | pes_2_13_io_stateOut == 4'h6 |
    pes_2_14_io_stateOut == 4'h6 | _T_159; // @[PEArray.scala 103:70]
  wire  _T_220 = pes_0_0_io_peconfig_ready | pes_0_1_io_peconfig_ready | pes_0_2_io_peconfig_ready |
    pes_0_3_io_peconfig_ready | pes_0_4_io_peconfig_ready | pes_0_5_io_peconfig_ready | pes_0_6_io_peconfig_ready |
    pes_0_7_io_peconfig_ready | pes_0_8_io_peconfig_ready | pes_0_9_io_peconfig_ready | pes_0_10_io_peconfig_ready |
    pes_0_11_io_peconfig_ready | pes_0_12_io_peconfig_ready | pes_0_13_io_peconfig_ready | pes_0_14_io_peconfig_ready |
    pes_0_15_io_peconfig_ready | pes_0_16_io_peconfig_ready | pes_0_17_io_peconfig_ready | pes_0_18_io_peconfig_ready |
    pes_0_19_io_peconfig_ready | pes_0_20_io_peconfig_ready | pes_0_21_io_peconfig_ready | pes_0_22_io_peconfig_ready |
    pes_0_23_io_peconfig_ready | pes_1_0_io_peconfig_ready | pes_1_1_io_peconfig_ready | pes_1_2_io_peconfig_ready |
    pes_1_3_io_peconfig_ready | pes_1_4_io_peconfig_ready | pes_1_5_io_peconfig_ready | pes_1_6_io_peconfig_ready; // @[PEArray.scala 106:77]
  wire  _T_250 = _T_220 | pes_1_7_io_peconfig_ready | pes_1_8_io_peconfig_ready | pes_1_9_io_peconfig_ready |
    pes_1_10_io_peconfig_ready | pes_1_11_io_peconfig_ready | pes_1_12_io_peconfig_ready | pes_1_13_io_peconfig_ready |
    pes_1_14_io_peconfig_ready | pes_1_15_io_peconfig_ready | pes_1_16_io_peconfig_ready | pes_1_17_io_peconfig_ready |
    pes_1_18_io_peconfig_ready | pes_1_19_io_peconfig_ready | pes_1_20_io_peconfig_ready | pes_1_21_io_peconfig_ready |
    pes_1_22_io_peconfig_ready | pes_1_23_io_peconfig_ready | pes_2_0_io_peconfig_ready | pes_2_1_io_peconfig_ready |
    pes_2_2_io_peconfig_ready | pes_2_3_io_peconfig_ready | pes_2_4_io_peconfig_ready | pes_2_5_io_peconfig_ready |
    pes_2_6_io_peconfig_ready | pes_2_7_io_peconfig_ready | pes_2_8_io_peconfig_ready | pes_2_9_io_peconfig_ready |
    pes_2_10_io_peconfig_ready | pes_2_11_io_peconfig_ready | pes_2_12_io_peconfig_ready; // @[PEArray.scala 106:77]
  Node NoC_0_0 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_0_clock),
    .reset(NoC_0_0_reset),
    .io_dataPackageIn_ready(NoC_0_0_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_0_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_0_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_0_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_row(NoC_0_0_io_dataPackageIn_bits_positon_row),
    .io_dataPackageIn_bits_positon_col(NoC_0_0_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_0_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_0_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_0_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_0_io_dataPackageOut_bits_dataType),
    .io_dataPackageOut_bits_positon_col(NoC_0_0_io_dataPackageOut_bits_positon_col)
  );
  Node_1 NoC_0_1 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_1_clock),
    .reset(NoC_0_1_reset),
    .io_dataPackageIn_ready(NoC_0_1_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_1_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_1_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_1_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_1_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_1_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_1_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_1_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_1_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_0 ( // @[PEArray.scala 36:24]
    .clock(pes_0_0_clock),
    .reset(pes_0_0_reset),
    .io_stateSW(pes_0_0_io_stateSW),
    .io_peconfig_ready(pes_0_0_io_peconfig_ready),
    .io_peconfig_valid(pes_0_0_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_0_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_0_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_0_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_0_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_0_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_0_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_0_io_filter_ready),
    .io_filter_valid(pes_0_0_io_filter_valid),
    .io_filter_bits(pes_0_0_io_filter_bits),
    .io_ifmap_ready(pes_0_0_io_ifmap_ready),
    .io_ifmap_valid(pes_0_0_io_ifmap_valid),
    .io_ifmap_bits(pes_0_0_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_0_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_0_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_0_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_0_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_0_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_0_io_pSumOut_bits),
    .io_stateOut(pes_0_0_io_stateOut)
  );
  dataSwitch dss_0_0 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_0_io_dataIn_ready),
    .io_dataIn_valid(dss_0_0_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_0_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_0_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_0_io_filter_ready),
    .io_filter_valid(dss_0_0_io_filter_valid),
    .io_filter_bits(dss_0_0_io_filter_bits),
    .io_ifmap_ready(dss_0_0_io_ifmap_ready),
    .io_ifmap_valid(dss_0_0_io_ifmap_valid),
    .io_ifmap_bits(dss_0_0_io_ifmap_bits),
    .io_pSum_ready(dss_0_0_io_pSum_ready),
    .io_pSum_valid(dss_0_0_io_pSum_valid),
    .io_pSum_bits(dss_0_0_io_pSum_bits)
  );
  Node_2 NoC_0_2 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_2_clock),
    .reset(NoC_0_2_reset),
    .io_dataPackageIn_ready(NoC_0_2_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_2_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_2_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_2_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_2_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_2_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_2_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_2_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_2_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_1 ( // @[PEArray.scala 36:24]
    .clock(pes_0_1_clock),
    .reset(pes_0_1_reset),
    .io_stateSW(pes_0_1_io_stateSW),
    .io_peconfig_ready(pes_0_1_io_peconfig_ready),
    .io_peconfig_valid(pes_0_1_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_1_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_1_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_1_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_1_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_1_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_1_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_1_io_filter_ready),
    .io_filter_valid(pes_0_1_io_filter_valid),
    .io_filter_bits(pes_0_1_io_filter_bits),
    .io_ifmap_ready(pes_0_1_io_ifmap_ready),
    .io_ifmap_valid(pes_0_1_io_ifmap_valid),
    .io_ifmap_bits(pes_0_1_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_1_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_1_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_1_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_1_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_1_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_1_io_pSumOut_bits),
    .io_stateOut(pes_0_1_io_stateOut)
  );
  dataSwitch dss_0_1 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_1_io_dataIn_ready),
    .io_dataIn_valid(dss_0_1_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_1_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_1_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_1_io_filter_ready),
    .io_filter_valid(dss_0_1_io_filter_valid),
    .io_filter_bits(dss_0_1_io_filter_bits),
    .io_ifmap_ready(dss_0_1_io_ifmap_ready),
    .io_ifmap_valid(dss_0_1_io_ifmap_valid),
    .io_ifmap_bits(dss_0_1_io_ifmap_bits),
    .io_pSum_ready(dss_0_1_io_pSum_ready),
    .io_pSum_valid(dss_0_1_io_pSum_valid),
    .io_pSum_bits(dss_0_1_io_pSum_bits)
  );
  Node_3 NoC_0_3 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_3_clock),
    .reset(NoC_0_3_reset),
    .io_dataPackageIn_ready(NoC_0_3_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_3_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_3_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_3_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_3_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_3_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_3_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_3_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_3_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_2 ( // @[PEArray.scala 36:24]
    .clock(pes_0_2_clock),
    .reset(pes_0_2_reset),
    .io_stateSW(pes_0_2_io_stateSW),
    .io_peconfig_ready(pes_0_2_io_peconfig_ready),
    .io_peconfig_valid(pes_0_2_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_2_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_2_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_2_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_2_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_2_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_2_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_2_io_filter_ready),
    .io_filter_valid(pes_0_2_io_filter_valid),
    .io_filter_bits(pes_0_2_io_filter_bits),
    .io_ifmap_ready(pes_0_2_io_ifmap_ready),
    .io_ifmap_valid(pes_0_2_io_ifmap_valid),
    .io_ifmap_bits(pes_0_2_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_2_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_2_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_2_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_2_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_2_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_2_io_pSumOut_bits),
    .io_stateOut(pes_0_2_io_stateOut)
  );
  dataSwitch dss_0_2 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_2_io_dataIn_ready),
    .io_dataIn_valid(dss_0_2_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_2_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_2_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_2_io_filter_ready),
    .io_filter_valid(dss_0_2_io_filter_valid),
    .io_filter_bits(dss_0_2_io_filter_bits),
    .io_ifmap_ready(dss_0_2_io_ifmap_ready),
    .io_ifmap_valid(dss_0_2_io_ifmap_valid),
    .io_ifmap_bits(dss_0_2_io_ifmap_bits),
    .io_pSum_ready(dss_0_2_io_pSum_ready),
    .io_pSum_valid(dss_0_2_io_pSum_valid),
    .io_pSum_bits(dss_0_2_io_pSum_bits)
  );
  Node_4 NoC_0_4 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_4_clock),
    .reset(NoC_0_4_reset),
    .io_dataPackageIn_ready(NoC_0_4_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_4_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_4_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_4_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_4_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_4_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_4_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_4_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_4_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_3 ( // @[PEArray.scala 36:24]
    .clock(pes_0_3_clock),
    .reset(pes_0_3_reset),
    .io_stateSW(pes_0_3_io_stateSW),
    .io_peconfig_ready(pes_0_3_io_peconfig_ready),
    .io_peconfig_valid(pes_0_3_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_3_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_3_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_3_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_3_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_3_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_3_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_3_io_filter_ready),
    .io_filter_valid(pes_0_3_io_filter_valid),
    .io_filter_bits(pes_0_3_io_filter_bits),
    .io_ifmap_ready(pes_0_3_io_ifmap_ready),
    .io_ifmap_valid(pes_0_3_io_ifmap_valid),
    .io_ifmap_bits(pes_0_3_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_3_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_3_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_3_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_3_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_3_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_3_io_pSumOut_bits),
    .io_stateOut(pes_0_3_io_stateOut)
  );
  dataSwitch dss_0_3 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_3_io_dataIn_ready),
    .io_dataIn_valid(dss_0_3_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_3_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_3_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_3_io_filter_ready),
    .io_filter_valid(dss_0_3_io_filter_valid),
    .io_filter_bits(dss_0_3_io_filter_bits),
    .io_ifmap_ready(dss_0_3_io_ifmap_ready),
    .io_ifmap_valid(dss_0_3_io_ifmap_valid),
    .io_ifmap_bits(dss_0_3_io_ifmap_bits),
    .io_pSum_ready(dss_0_3_io_pSum_ready),
    .io_pSum_valid(dss_0_3_io_pSum_valid),
    .io_pSum_bits(dss_0_3_io_pSum_bits)
  );
  Node_5 NoC_0_5 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_5_clock),
    .reset(NoC_0_5_reset),
    .io_dataPackageIn_ready(NoC_0_5_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_5_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_5_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_5_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_5_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_5_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_5_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_5_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_5_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_4 ( // @[PEArray.scala 36:24]
    .clock(pes_0_4_clock),
    .reset(pes_0_4_reset),
    .io_stateSW(pes_0_4_io_stateSW),
    .io_peconfig_ready(pes_0_4_io_peconfig_ready),
    .io_peconfig_valid(pes_0_4_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_4_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_4_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_4_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_4_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_4_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_4_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_4_io_filter_ready),
    .io_filter_valid(pes_0_4_io_filter_valid),
    .io_filter_bits(pes_0_4_io_filter_bits),
    .io_ifmap_ready(pes_0_4_io_ifmap_ready),
    .io_ifmap_valid(pes_0_4_io_ifmap_valid),
    .io_ifmap_bits(pes_0_4_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_4_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_4_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_4_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_4_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_4_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_4_io_pSumOut_bits),
    .io_stateOut(pes_0_4_io_stateOut)
  );
  dataSwitch dss_0_4 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_4_io_dataIn_ready),
    .io_dataIn_valid(dss_0_4_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_4_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_4_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_4_io_filter_ready),
    .io_filter_valid(dss_0_4_io_filter_valid),
    .io_filter_bits(dss_0_4_io_filter_bits),
    .io_ifmap_ready(dss_0_4_io_ifmap_ready),
    .io_ifmap_valid(dss_0_4_io_ifmap_valid),
    .io_ifmap_bits(dss_0_4_io_ifmap_bits),
    .io_pSum_ready(dss_0_4_io_pSum_ready),
    .io_pSum_valid(dss_0_4_io_pSum_valid),
    .io_pSum_bits(dss_0_4_io_pSum_bits)
  );
  Node_6 NoC_0_6 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_6_clock),
    .reset(NoC_0_6_reset),
    .io_dataPackageIn_ready(NoC_0_6_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_6_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_6_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_6_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_6_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_6_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_6_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_6_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_6_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_5 ( // @[PEArray.scala 36:24]
    .clock(pes_0_5_clock),
    .reset(pes_0_5_reset),
    .io_stateSW(pes_0_5_io_stateSW),
    .io_peconfig_ready(pes_0_5_io_peconfig_ready),
    .io_peconfig_valid(pes_0_5_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_5_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_5_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_5_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_5_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_5_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_5_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_5_io_filter_ready),
    .io_filter_valid(pes_0_5_io_filter_valid),
    .io_filter_bits(pes_0_5_io_filter_bits),
    .io_ifmap_ready(pes_0_5_io_ifmap_ready),
    .io_ifmap_valid(pes_0_5_io_ifmap_valid),
    .io_ifmap_bits(pes_0_5_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_5_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_5_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_5_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_5_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_5_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_5_io_pSumOut_bits),
    .io_stateOut(pes_0_5_io_stateOut)
  );
  dataSwitch dss_0_5 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_5_io_dataIn_ready),
    .io_dataIn_valid(dss_0_5_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_5_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_5_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_5_io_filter_ready),
    .io_filter_valid(dss_0_5_io_filter_valid),
    .io_filter_bits(dss_0_5_io_filter_bits),
    .io_ifmap_ready(dss_0_5_io_ifmap_ready),
    .io_ifmap_valid(dss_0_5_io_ifmap_valid),
    .io_ifmap_bits(dss_0_5_io_ifmap_bits),
    .io_pSum_ready(dss_0_5_io_pSum_ready),
    .io_pSum_valid(dss_0_5_io_pSum_valid),
    .io_pSum_bits(dss_0_5_io_pSum_bits)
  );
  Node_7 NoC_0_7 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_7_clock),
    .reset(NoC_0_7_reset),
    .io_dataPackageIn_ready(NoC_0_7_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_7_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_7_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_7_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_7_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_7_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_7_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_7_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_7_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_6 ( // @[PEArray.scala 36:24]
    .clock(pes_0_6_clock),
    .reset(pes_0_6_reset),
    .io_stateSW(pes_0_6_io_stateSW),
    .io_peconfig_ready(pes_0_6_io_peconfig_ready),
    .io_peconfig_valid(pes_0_6_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_6_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_6_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_6_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_6_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_6_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_6_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_6_io_filter_ready),
    .io_filter_valid(pes_0_6_io_filter_valid),
    .io_filter_bits(pes_0_6_io_filter_bits),
    .io_ifmap_ready(pes_0_6_io_ifmap_ready),
    .io_ifmap_valid(pes_0_6_io_ifmap_valid),
    .io_ifmap_bits(pes_0_6_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_6_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_6_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_6_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_6_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_6_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_6_io_pSumOut_bits),
    .io_stateOut(pes_0_6_io_stateOut)
  );
  dataSwitch dss_0_6 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_6_io_dataIn_ready),
    .io_dataIn_valid(dss_0_6_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_6_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_6_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_6_io_filter_ready),
    .io_filter_valid(dss_0_6_io_filter_valid),
    .io_filter_bits(dss_0_6_io_filter_bits),
    .io_ifmap_ready(dss_0_6_io_ifmap_ready),
    .io_ifmap_valid(dss_0_6_io_ifmap_valid),
    .io_ifmap_bits(dss_0_6_io_ifmap_bits),
    .io_pSum_ready(dss_0_6_io_pSum_ready),
    .io_pSum_valid(dss_0_6_io_pSum_valid),
    .io_pSum_bits(dss_0_6_io_pSum_bits)
  );
  Node_8 NoC_0_8 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_8_clock),
    .reset(NoC_0_8_reset),
    .io_dataPackageIn_ready(NoC_0_8_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_8_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_8_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_8_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_8_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_8_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_8_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_8_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_8_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_7 ( // @[PEArray.scala 36:24]
    .clock(pes_0_7_clock),
    .reset(pes_0_7_reset),
    .io_stateSW(pes_0_7_io_stateSW),
    .io_peconfig_ready(pes_0_7_io_peconfig_ready),
    .io_peconfig_valid(pes_0_7_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_7_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_7_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_7_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_7_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_7_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_7_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_7_io_filter_ready),
    .io_filter_valid(pes_0_7_io_filter_valid),
    .io_filter_bits(pes_0_7_io_filter_bits),
    .io_ifmap_ready(pes_0_7_io_ifmap_ready),
    .io_ifmap_valid(pes_0_7_io_ifmap_valid),
    .io_ifmap_bits(pes_0_7_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_7_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_7_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_7_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_7_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_7_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_7_io_pSumOut_bits),
    .io_stateOut(pes_0_7_io_stateOut)
  );
  dataSwitch dss_0_7 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_7_io_dataIn_ready),
    .io_dataIn_valid(dss_0_7_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_7_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_7_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_7_io_filter_ready),
    .io_filter_valid(dss_0_7_io_filter_valid),
    .io_filter_bits(dss_0_7_io_filter_bits),
    .io_ifmap_ready(dss_0_7_io_ifmap_ready),
    .io_ifmap_valid(dss_0_7_io_ifmap_valid),
    .io_ifmap_bits(dss_0_7_io_ifmap_bits),
    .io_pSum_ready(dss_0_7_io_pSum_ready),
    .io_pSum_valid(dss_0_7_io_pSum_valid),
    .io_pSum_bits(dss_0_7_io_pSum_bits)
  );
  Node_9 NoC_0_9 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_9_clock),
    .reset(NoC_0_9_reset),
    .io_dataPackageIn_ready(NoC_0_9_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_9_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_9_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_9_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_9_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_9_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_9_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_9_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_9_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_8 ( // @[PEArray.scala 36:24]
    .clock(pes_0_8_clock),
    .reset(pes_0_8_reset),
    .io_stateSW(pes_0_8_io_stateSW),
    .io_peconfig_ready(pes_0_8_io_peconfig_ready),
    .io_peconfig_valid(pes_0_8_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_8_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_8_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_8_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_8_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_8_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_8_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_8_io_filter_ready),
    .io_filter_valid(pes_0_8_io_filter_valid),
    .io_filter_bits(pes_0_8_io_filter_bits),
    .io_ifmap_ready(pes_0_8_io_ifmap_ready),
    .io_ifmap_valid(pes_0_8_io_ifmap_valid),
    .io_ifmap_bits(pes_0_8_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_8_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_8_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_8_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_8_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_8_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_8_io_pSumOut_bits),
    .io_stateOut(pes_0_8_io_stateOut)
  );
  dataSwitch dss_0_8 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_8_io_dataIn_ready),
    .io_dataIn_valid(dss_0_8_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_8_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_8_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_8_io_filter_ready),
    .io_filter_valid(dss_0_8_io_filter_valid),
    .io_filter_bits(dss_0_8_io_filter_bits),
    .io_ifmap_ready(dss_0_8_io_ifmap_ready),
    .io_ifmap_valid(dss_0_8_io_ifmap_valid),
    .io_ifmap_bits(dss_0_8_io_ifmap_bits),
    .io_pSum_ready(dss_0_8_io_pSum_ready),
    .io_pSum_valid(dss_0_8_io_pSum_valid),
    .io_pSum_bits(dss_0_8_io_pSum_bits)
  );
  Node_10 NoC_0_10 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_10_clock),
    .reset(NoC_0_10_reset),
    .io_dataPackageIn_ready(NoC_0_10_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_10_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_10_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_10_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_10_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_10_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_10_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_10_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_10_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_9 ( // @[PEArray.scala 36:24]
    .clock(pes_0_9_clock),
    .reset(pes_0_9_reset),
    .io_stateSW(pes_0_9_io_stateSW),
    .io_peconfig_ready(pes_0_9_io_peconfig_ready),
    .io_peconfig_valid(pes_0_9_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_9_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_9_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_9_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_9_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_9_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_9_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_9_io_filter_ready),
    .io_filter_valid(pes_0_9_io_filter_valid),
    .io_filter_bits(pes_0_9_io_filter_bits),
    .io_ifmap_ready(pes_0_9_io_ifmap_ready),
    .io_ifmap_valid(pes_0_9_io_ifmap_valid),
    .io_ifmap_bits(pes_0_9_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_9_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_9_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_9_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_9_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_9_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_9_io_pSumOut_bits),
    .io_stateOut(pes_0_9_io_stateOut)
  );
  dataSwitch dss_0_9 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_9_io_dataIn_ready),
    .io_dataIn_valid(dss_0_9_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_9_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_9_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_9_io_filter_ready),
    .io_filter_valid(dss_0_9_io_filter_valid),
    .io_filter_bits(dss_0_9_io_filter_bits),
    .io_ifmap_ready(dss_0_9_io_ifmap_ready),
    .io_ifmap_valid(dss_0_9_io_ifmap_valid),
    .io_ifmap_bits(dss_0_9_io_ifmap_bits),
    .io_pSum_ready(dss_0_9_io_pSum_ready),
    .io_pSum_valid(dss_0_9_io_pSum_valid),
    .io_pSum_bits(dss_0_9_io_pSum_bits)
  );
  Node_11 NoC_0_11 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_11_clock),
    .reset(NoC_0_11_reset),
    .io_dataPackageIn_ready(NoC_0_11_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_11_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_11_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_11_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_11_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_11_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_11_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_11_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_11_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_10 ( // @[PEArray.scala 36:24]
    .clock(pes_0_10_clock),
    .reset(pes_0_10_reset),
    .io_stateSW(pes_0_10_io_stateSW),
    .io_peconfig_ready(pes_0_10_io_peconfig_ready),
    .io_peconfig_valid(pes_0_10_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_10_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_10_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_10_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_10_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_10_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_10_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_10_io_filter_ready),
    .io_filter_valid(pes_0_10_io_filter_valid),
    .io_filter_bits(pes_0_10_io_filter_bits),
    .io_ifmap_ready(pes_0_10_io_ifmap_ready),
    .io_ifmap_valid(pes_0_10_io_ifmap_valid),
    .io_ifmap_bits(pes_0_10_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_10_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_10_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_10_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_10_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_10_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_10_io_pSumOut_bits),
    .io_stateOut(pes_0_10_io_stateOut)
  );
  dataSwitch dss_0_10 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_10_io_dataIn_ready),
    .io_dataIn_valid(dss_0_10_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_10_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_10_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_10_io_filter_ready),
    .io_filter_valid(dss_0_10_io_filter_valid),
    .io_filter_bits(dss_0_10_io_filter_bits),
    .io_ifmap_ready(dss_0_10_io_ifmap_ready),
    .io_ifmap_valid(dss_0_10_io_ifmap_valid),
    .io_ifmap_bits(dss_0_10_io_ifmap_bits),
    .io_pSum_ready(dss_0_10_io_pSum_ready),
    .io_pSum_valid(dss_0_10_io_pSum_valid),
    .io_pSum_bits(dss_0_10_io_pSum_bits)
  );
  Node_12 NoC_0_12 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_12_clock),
    .reset(NoC_0_12_reset),
    .io_dataPackageIn_ready(NoC_0_12_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_12_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_12_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_12_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_12_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_12_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_12_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_12_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_12_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_11 ( // @[PEArray.scala 36:24]
    .clock(pes_0_11_clock),
    .reset(pes_0_11_reset),
    .io_stateSW(pes_0_11_io_stateSW),
    .io_peconfig_ready(pes_0_11_io_peconfig_ready),
    .io_peconfig_valid(pes_0_11_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_11_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_11_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_11_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_11_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_11_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_11_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_11_io_filter_ready),
    .io_filter_valid(pes_0_11_io_filter_valid),
    .io_filter_bits(pes_0_11_io_filter_bits),
    .io_ifmap_ready(pes_0_11_io_ifmap_ready),
    .io_ifmap_valid(pes_0_11_io_ifmap_valid),
    .io_ifmap_bits(pes_0_11_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_11_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_11_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_11_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_11_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_11_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_11_io_pSumOut_bits),
    .io_stateOut(pes_0_11_io_stateOut)
  );
  dataSwitch dss_0_11 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_11_io_dataIn_ready),
    .io_dataIn_valid(dss_0_11_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_11_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_11_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_11_io_filter_ready),
    .io_filter_valid(dss_0_11_io_filter_valid),
    .io_filter_bits(dss_0_11_io_filter_bits),
    .io_ifmap_ready(dss_0_11_io_ifmap_ready),
    .io_ifmap_valid(dss_0_11_io_ifmap_valid),
    .io_ifmap_bits(dss_0_11_io_ifmap_bits),
    .io_pSum_ready(dss_0_11_io_pSum_ready),
    .io_pSum_valid(dss_0_11_io_pSum_valid),
    .io_pSum_bits(dss_0_11_io_pSum_bits)
  );
  Node_13 NoC_0_13 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_13_clock),
    .reset(NoC_0_13_reset),
    .io_dataPackageIn_ready(NoC_0_13_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_13_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_13_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_13_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_13_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_13_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_13_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_13_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_13_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_12 ( // @[PEArray.scala 36:24]
    .clock(pes_0_12_clock),
    .reset(pes_0_12_reset),
    .io_stateSW(pes_0_12_io_stateSW),
    .io_peconfig_ready(pes_0_12_io_peconfig_ready),
    .io_peconfig_valid(pes_0_12_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_12_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_12_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_12_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_12_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_12_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_12_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_12_io_filter_ready),
    .io_filter_valid(pes_0_12_io_filter_valid),
    .io_filter_bits(pes_0_12_io_filter_bits),
    .io_ifmap_ready(pes_0_12_io_ifmap_ready),
    .io_ifmap_valid(pes_0_12_io_ifmap_valid),
    .io_ifmap_bits(pes_0_12_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_12_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_12_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_12_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_12_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_12_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_12_io_pSumOut_bits),
    .io_stateOut(pes_0_12_io_stateOut)
  );
  dataSwitch dss_0_12 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_12_io_dataIn_ready),
    .io_dataIn_valid(dss_0_12_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_12_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_12_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_12_io_filter_ready),
    .io_filter_valid(dss_0_12_io_filter_valid),
    .io_filter_bits(dss_0_12_io_filter_bits),
    .io_ifmap_ready(dss_0_12_io_ifmap_ready),
    .io_ifmap_valid(dss_0_12_io_ifmap_valid),
    .io_ifmap_bits(dss_0_12_io_ifmap_bits),
    .io_pSum_ready(dss_0_12_io_pSum_ready),
    .io_pSum_valid(dss_0_12_io_pSum_valid),
    .io_pSum_bits(dss_0_12_io_pSum_bits)
  );
  Node_14 NoC_0_14 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_14_clock),
    .reset(NoC_0_14_reset),
    .io_dataPackageIn_ready(NoC_0_14_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_14_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_14_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_14_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_14_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_14_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_14_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_14_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_14_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_13 ( // @[PEArray.scala 36:24]
    .clock(pes_0_13_clock),
    .reset(pes_0_13_reset),
    .io_stateSW(pes_0_13_io_stateSW),
    .io_peconfig_ready(pes_0_13_io_peconfig_ready),
    .io_peconfig_valid(pes_0_13_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_13_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_13_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_13_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_13_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_13_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_13_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_13_io_filter_ready),
    .io_filter_valid(pes_0_13_io_filter_valid),
    .io_filter_bits(pes_0_13_io_filter_bits),
    .io_ifmap_ready(pes_0_13_io_ifmap_ready),
    .io_ifmap_valid(pes_0_13_io_ifmap_valid),
    .io_ifmap_bits(pes_0_13_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_13_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_13_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_13_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_13_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_13_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_13_io_pSumOut_bits),
    .io_stateOut(pes_0_13_io_stateOut)
  );
  dataSwitch dss_0_13 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_13_io_dataIn_ready),
    .io_dataIn_valid(dss_0_13_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_13_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_13_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_13_io_filter_ready),
    .io_filter_valid(dss_0_13_io_filter_valid),
    .io_filter_bits(dss_0_13_io_filter_bits),
    .io_ifmap_ready(dss_0_13_io_ifmap_ready),
    .io_ifmap_valid(dss_0_13_io_ifmap_valid),
    .io_ifmap_bits(dss_0_13_io_ifmap_bits),
    .io_pSum_ready(dss_0_13_io_pSum_ready),
    .io_pSum_valid(dss_0_13_io_pSum_valid),
    .io_pSum_bits(dss_0_13_io_pSum_bits)
  );
  Node_15 NoC_0_15 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_15_clock),
    .reset(NoC_0_15_reset),
    .io_dataPackageIn_ready(NoC_0_15_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_15_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_15_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_15_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_15_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_15_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_15_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_15_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_15_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_14 ( // @[PEArray.scala 36:24]
    .clock(pes_0_14_clock),
    .reset(pes_0_14_reset),
    .io_stateSW(pes_0_14_io_stateSW),
    .io_peconfig_ready(pes_0_14_io_peconfig_ready),
    .io_peconfig_valid(pes_0_14_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_14_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_14_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_14_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_14_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_14_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_14_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_14_io_filter_ready),
    .io_filter_valid(pes_0_14_io_filter_valid),
    .io_filter_bits(pes_0_14_io_filter_bits),
    .io_ifmap_ready(pes_0_14_io_ifmap_ready),
    .io_ifmap_valid(pes_0_14_io_ifmap_valid),
    .io_ifmap_bits(pes_0_14_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_14_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_14_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_14_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_14_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_14_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_14_io_pSumOut_bits),
    .io_stateOut(pes_0_14_io_stateOut)
  );
  dataSwitch dss_0_14 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_14_io_dataIn_ready),
    .io_dataIn_valid(dss_0_14_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_14_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_14_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_14_io_filter_ready),
    .io_filter_valid(dss_0_14_io_filter_valid),
    .io_filter_bits(dss_0_14_io_filter_bits),
    .io_ifmap_ready(dss_0_14_io_ifmap_ready),
    .io_ifmap_valid(dss_0_14_io_ifmap_valid),
    .io_ifmap_bits(dss_0_14_io_ifmap_bits),
    .io_pSum_ready(dss_0_14_io_pSum_ready),
    .io_pSum_valid(dss_0_14_io_pSum_valid),
    .io_pSum_bits(dss_0_14_io_pSum_bits)
  );
  Node_16 NoC_0_16 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_16_clock),
    .reset(NoC_0_16_reset),
    .io_dataPackageIn_ready(NoC_0_16_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_16_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_16_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_16_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_16_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_16_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_16_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_16_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_16_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_15 ( // @[PEArray.scala 36:24]
    .clock(pes_0_15_clock),
    .reset(pes_0_15_reset),
    .io_stateSW(pes_0_15_io_stateSW),
    .io_peconfig_ready(pes_0_15_io_peconfig_ready),
    .io_peconfig_valid(pes_0_15_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_15_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_15_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_15_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_15_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_15_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_15_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_15_io_filter_ready),
    .io_filter_valid(pes_0_15_io_filter_valid),
    .io_filter_bits(pes_0_15_io_filter_bits),
    .io_ifmap_ready(pes_0_15_io_ifmap_ready),
    .io_ifmap_valid(pes_0_15_io_ifmap_valid),
    .io_ifmap_bits(pes_0_15_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_15_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_15_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_15_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_15_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_15_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_15_io_pSumOut_bits),
    .io_stateOut(pes_0_15_io_stateOut)
  );
  dataSwitch dss_0_15 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_15_io_dataIn_ready),
    .io_dataIn_valid(dss_0_15_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_15_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_15_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_15_io_filter_ready),
    .io_filter_valid(dss_0_15_io_filter_valid),
    .io_filter_bits(dss_0_15_io_filter_bits),
    .io_ifmap_ready(dss_0_15_io_ifmap_ready),
    .io_ifmap_valid(dss_0_15_io_ifmap_valid),
    .io_ifmap_bits(dss_0_15_io_ifmap_bits),
    .io_pSum_ready(dss_0_15_io_pSum_ready),
    .io_pSum_valid(dss_0_15_io_pSum_valid),
    .io_pSum_bits(dss_0_15_io_pSum_bits)
  );
  Node_17 NoC_0_17 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_17_clock),
    .reset(NoC_0_17_reset),
    .io_dataPackageIn_ready(NoC_0_17_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_17_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_17_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_17_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_17_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_17_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_17_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_17_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_17_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_16 ( // @[PEArray.scala 36:24]
    .clock(pes_0_16_clock),
    .reset(pes_0_16_reset),
    .io_stateSW(pes_0_16_io_stateSW),
    .io_peconfig_ready(pes_0_16_io_peconfig_ready),
    .io_peconfig_valid(pes_0_16_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_16_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_16_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_16_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_16_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_16_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_16_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_16_io_filter_ready),
    .io_filter_valid(pes_0_16_io_filter_valid),
    .io_filter_bits(pes_0_16_io_filter_bits),
    .io_ifmap_ready(pes_0_16_io_ifmap_ready),
    .io_ifmap_valid(pes_0_16_io_ifmap_valid),
    .io_ifmap_bits(pes_0_16_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_16_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_16_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_16_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_16_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_16_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_16_io_pSumOut_bits),
    .io_stateOut(pes_0_16_io_stateOut)
  );
  dataSwitch dss_0_16 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_16_io_dataIn_ready),
    .io_dataIn_valid(dss_0_16_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_16_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_16_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_16_io_filter_ready),
    .io_filter_valid(dss_0_16_io_filter_valid),
    .io_filter_bits(dss_0_16_io_filter_bits),
    .io_ifmap_ready(dss_0_16_io_ifmap_ready),
    .io_ifmap_valid(dss_0_16_io_ifmap_valid),
    .io_ifmap_bits(dss_0_16_io_ifmap_bits),
    .io_pSum_ready(dss_0_16_io_pSum_ready),
    .io_pSum_valid(dss_0_16_io_pSum_valid),
    .io_pSum_bits(dss_0_16_io_pSum_bits)
  );
  Node_18 NoC_0_18 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_18_clock),
    .reset(NoC_0_18_reset),
    .io_dataPackageIn_ready(NoC_0_18_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_18_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_18_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_18_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_18_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_18_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_18_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_18_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_18_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_17 ( // @[PEArray.scala 36:24]
    .clock(pes_0_17_clock),
    .reset(pes_0_17_reset),
    .io_stateSW(pes_0_17_io_stateSW),
    .io_peconfig_ready(pes_0_17_io_peconfig_ready),
    .io_peconfig_valid(pes_0_17_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_17_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_17_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_17_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_17_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_17_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_17_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_17_io_filter_ready),
    .io_filter_valid(pes_0_17_io_filter_valid),
    .io_filter_bits(pes_0_17_io_filter_bits),
    .io_ifmap_ready(pes_0_17_io_ifmap_ready),
    .io_ifmap_valid(pes_0_17_io_ifmap_valid),
    .io_ifmap_bits(pes_0_17_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_17_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_17_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_17_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_17_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_17_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_17_io_pSumOut_bits),
    .io_stateOut(pes_0_17_io_stateOut)
  );
  dataSwitch dss_0_17 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_17_io_dataIn_ready),
    .io_dataIn_valid(dss_0_17_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_17_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_17_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_17_io_filter_ready),
    .io_filter_valid(dss_0_17_io_filter_valid),
    .io_filter_bits(dss_0_17_io_filter_bits),
    .io_ifmap_ready(dss_0_17_io_ifmap_ready),
    .io_ifmap_valid(dss_0_17_io_ifmap_valid),
    .io_ifmap_bits(dss_0_17_io_ifmap_bits),
    .io_pSum_ready(dss_0_17_io_pSum_ready),
    .io_pSum_valid(dss_0_17_io_pSum_valid),
    .io_pSum_bits(dss_0_17_io_pSum_bits)
  );
  Node_19 NoC_0_19 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_19_clock),
    .reset(NoC_0_19_reset),
    .io_dataPackageIn_ready(NoC_0_19_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_19_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_19_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_19_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_19_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_19_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_19_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_19_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_19_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_18 ( // @[PEArray.scala 36:24]
    .clock(pes_0_18_clock),
    .reset(pes_0_18_reset),
    .io_stateSW(pes_0_18_io_stateSW),
    .io_peconfig_ready(pes_0_18_io_peconfig_ready),
    .io_peconfig_valid(pes_0_18_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_18_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_18_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_18_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_18_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_18_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_18_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_18_io_filter_ready),
    .io_filter_valid(pes_0_18_io_filter_valid),
    .io_filter_bits(pes_0_18_io_filter_bits),
    .io_ifmap_ready(pes_0_18_io_ifmap_ready),
    .io_ifmap_valid(pes_0_18_io_ifmap_valid),
    .io_ifmap_bits(pes_0_18_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_18_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_18_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_18_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_18_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_18_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_18_io_pSumOut_bits),
    .io_stateOut(pes_0_18_io_stateOut)
  );
  dataSwitch dss_0_18 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_18_io_dataIn_ready),
    .io_dataIn_valid(dss_0_18_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_18_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_18_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_18_io_filter_ready),
    .io_filter_valid(dss_0_18_io_filter_valid),
    .io_filter_bits(dss_0_18_io_filter_bits),
    .io_ifmap_ready(dss_0_18_io_ifmap_ready),
    .io_ifmap_valid(dss_0_18_io_ifmap_valid),
    .io_ifmap_bits(dss_0_18_io_ifmap_bits),
    .io_pSum_ready(dss_0_18_io_pSum_ready),
    .io_pSum_valid(dss_0_18_io_pSum_valid),
    .io_pSum_bits(dss_0_18_io_pSum_bits)
  );
  Node_20 NoC_0_20 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_20_clock),
    .reset(NoC_0_20_reset),
    .io_dataPackageIn_ready(NoC_0_20_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_20_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_20_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_20_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_20_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_20_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_20_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_20_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_20_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_19 ( // @[PEArray.scala 36:24]
    .clock(pes_0_19_clock),
    .reset(pes_0_19_reset),
    .io_stateSW(pes_0_19_io_stateSW),
    .io_peconfig_ready(pes_0_19_io_peconfig_ready),
    .io_peconfig_valid(pes_0_19_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_19_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_19_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_19_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_19_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_19_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_19_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_19_io_filter_ready),
    .io_filter_valid(pes_0_19_io_filter_valid),
    .io_filter_bits(pes_0_19_io_filter_bits),
    .io_ifmap_ready(pes_0_19_io_ifmap_ready),
    .io_ifmap_valid(pes_0_19_io_ifmap_valid),
    .io_ifmap_bits(pes_0_19_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_19_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_19_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_19_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_19_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_19_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_19_io_pSumOut_bits),
    .io_stateOut(pes_0_19_io_stateOut)
  );
  dataSwitch dss_0_19 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_19_io_dataIn_ready),
    .io_dataIn_valid(dss_0_19_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_19_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_19_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_19_io_filter_ready),
    .io_filter_valid(dss_0_19_io_filter_valid),
    .io_filter_bits(dss_0_19_io_filter_bits),
    .io_ifmap_ready(dss_0_19_io_ifmap_ready),
    .io_ifmap_valid(dss_0_19_io_ifmap_valid),
    .io_ifmap_bits(dss_0_19_io_ifmap_bits),
    .io_pSum_ready(dss_0_19_io_pSum_ready),
    .io_pSum_valid(dss_0_19_io_pSum_valid),
    .io_pSum_bits(dss_0_19_io_pSum_bits)
  );
  Node_21 NoC_0_21 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_21_clock),
    .reset(NoC_0_21_reset),
    .io_dataPackageIn_ready(NoC_0_21_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_21_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_21_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_21_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_21_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_21_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_21_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_21_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_21_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_20 ( // @[PEArray.scala 36:24]
    .clock(pes_0_20_clock),
    .reset(pes_0_20_reset),
    .io_stateSW(pes_0_20_io_stateSW),
    .io_peconfig_ready(pes_0_20_io_peconfig_ready),
    .io_peconfig_valid(pes_0_20_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_20_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_20_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_20_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_20_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_20_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_20_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_20_io_filter_ready),
    .io_filter_valid(pes_0_20_io_filter_valid),
    .io_filter_bits(pes_0_20_io_filter_bits),
    .io_ifmap_ready(pes_0_20_io_ifmap_ready),
    .io_ifmap_valid(pes_0_20_io_ifmap_valid),
    .io_ifmap_bits(pes_0_20_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_20_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_20_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_20_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_20_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_20_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_20_io_pSumOut_bits),
    .io_stateOut(pes_0_20_io_stateOut)
  );
  dataSwitch dss_0_20 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_20_io_dataIn_ready),
    .io_dataIn_valid(dss_0_20_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_20_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_20_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_20_io_filter_ready),
    .io_filter_valid(dss_0_20_io_filter_valid),
    .io_filter_bits(dss_0_20_io_filter_bits),
    .io_ifmap_ready(dss_0_20_io_ifmap_ready),
    .io_ifmap_valid(dss_0_20_io_ifmap_valid),
    .io_ifmap_bits(dss_0_20_io_ifmap_bits),
    .io_pSum_ready(dss_0_20_io_pSum_ready),
    .io_pSum_valid(dss_0_20_io_pSum_valid),
    .io_pSum_bits(dss_0_20_io_pSum_bits)
  );
  Node_22 NoC_0_22 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_22_clock),
    .reset(NoC_0_22_reset),
    .io_dataPackageIn_ready(NoC_0_22_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_22_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_22_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_22_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_22_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_22_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_22_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_22_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_22_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_21 ( // @[PEArray.scala 36:24]
    .clock(pes_0_21_clock),
    .reset(pes_0_21_reset),
    .io_stateSW(pes_0_21_io_stateSW),
    .io_peconfig_ready(pes_0_21_io_peconfig_ready),
    .io_peconfig_valid(pes_0_21_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_21_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_21_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_21_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_21_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_21_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_21_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_21_io_filter_ready),
    .io_filter_valid(pes_0_21_io_filter_valid),
    .io_filter_bits(pes_0_21_io_filter_bits),
    .io_ifmap_ready(pes_0_21_io_ifmap_ready),
    .io_ifmap_valid(pes_0_21_io_ifmap_valid),
    .io_ifmap_bits(pes_0_21_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_21_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_21_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_21_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_21_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_21_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_21_io_pSumOut_bits),
    .io_stateOut(pes_0_21_io_stateOut)
  );
  dataSwitch dss_0_21 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_21_io_dataIn_ready),
    .io_dataIn_valid(dss_0_21_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_21_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_21_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_21_io_filter_ready),
    .io_filter_valid(dss_0_21_io_filter_valid),
    .io_filter_bits(dss_0_21_io_filter_bits),
    .io_ifmap_ready(dss_0_21_io_ifmap_ready),
    .io_ifmap_valid(dss_0_21_io_ifmap_valid),
    .io_ifmap_bits(dss_0_21_io_ifmap_bits),
    .io_pSum_ready(dss_0_21_io_pSum_ready),
    .io_pSum_valid(dss_0_21_io_pSum_valid),
    .io_pSum_bits(dss_0_21_io_pSum_bits)
  );
  Node_23 NoC_0_23 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_23_clock),
    .reset(NoC_0_23_reset),
    .io_dataPackageIn_ready(NoC_0_23_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_23_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_23_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_23_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_23_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_23_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_23_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_23_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_23_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_22 ( // @[PEArray.scala 36:24]
    .clock(pes_0_22_clock),
    .reset(pes_0_22_reset),
    .io_stateSW(pes_0_22_io_stateSW),
    .io_peconfig_ready(pes_0_22_io_peconfig_ready),
    .io_peconfig_valid(pes_0_22_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_22_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_22_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_22_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_22_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_22_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_22_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_22_io_filter_ready),
    .io_filter_valid(pes_0_22_io_filter_valid),
    .io_filter_bits(pes_0_22_io_filter_bits),
    .io_ifmap_ready(pes_0_22_io_ifmap_ready),
    .io_ifmap_valid(pes_0_22_io_ifmap_valid),
    .io_ifmap_bits(pes_0_22_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_22_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_22_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_22_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_22_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_22_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_22_io_pSumOut_bits),
    .io_stateOut(pes_0_22_io_stateOut)
  );
  dataSwitch dss_0_22 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_22_io_dataIn_ready),
    .io_dataIn_valid(dss_0_22_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_22_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_22_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_22_io_filter_ready),
    .io_filter_valid(dss_0_22_io_filter_valid),
    .io_filter_bits(dss_0_22_io_filter_bits),
    .io_ifmap_ready(dss_0_22_io_ifmap_ready),
    .io_ifmap_valid(dss_0_22_io_ifmap_valid),
    .io_ifmap_bits(dss_0_22_io_ifmap_bits),
    .io_pSum_ready(dss_0_22_io_pSum_ready),
    .io_pSum_valid(dss_0_22_io_pSum_valid),
    .io_pSum_bits(dss_0_22_io_pSum_bits)
  );
  Node_24 NoC_0_24 ( // @[PEArray.scala 34:24]
    .clock(NoC_0_24_clock),
    .reset(NoC_0_24_reset),
    .io_dataPackageIn_ready(NoC_0_24_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_0_24_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_0_24_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_0_24_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_0_24_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_0_24_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_0_24_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_0_24_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_0_24_io_dataPackageOut_bits_dataType)
  );
  PETop pes_0_23 ( // @[PEArray.scala 36:24]
    .clock(pes_0_23_clock),
    .reset(pes_0_23_reset),
    .io_stateSW(pes_0_23_io_stateSW),
    .io_peconfig_ready(pes_0_23_io_peconfig_ready),
    .io_peconfig_valid(pes_0_23_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_0_23_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_0_23_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_0_23_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_0_23_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_0_23_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_0_23_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_0_23_io_filter_ready),
    .io_filter_valid(pes_0_23_io_filter_valid),
    .io_filter_bits(pes_0_23_io_filter_bits),
    .io_ifmap_ready(pes_0_23_io_ifmap_ready),
    .io_ifmap_valid(pes_0_23_io_ifmap_valid),
    .io_ifmap_bits(pes_0_23_io_ifmap_bits),
    .io_pSumIn_ready(pes_0_23_io_pSumIn_ready),
    .io_pSumIn_valid(pes_0_23_io_pSumIn_valid),
    .io_pSumIn_bits(pes_0_23_io_pSumIn_bits),
    .io_pSumOut_ready(pes_0_23_io_pSumOut_ready),
    .io_pSumOut_valid(pes_0_23_io_pSumOut_valid),
    .io_pSumOut_bits(pes_0_23_io_pSumOut_bits),
    .io_stateOut(pes_0_23_io_stateOut)
  );
  dataSwitch dss_0_23 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_0_23_io_dataIn_ready),
    .io_dataIn_valid(dss_0_23_io_dataIn_valid),
    .io_dataIn_bits_data(dss_0_23_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_0_23_io_dataIn_bits_dataType),
    .io_filter_ready(dss_0_23_io_filter_ready),
    .io_filter_valid(dss_0_23_io_filter_valid),
    .io_filter_bits(dss_0_23_io_filter_bits),
    .io_ifmap_ready(dss_0_23_io_ifmap_ready),
    .io_ifmap_valid(dss_0_23_io_ifmap_valid),
    .io_ifmap_bits(dss_0_23_io_ifmap_bits),
    .io_pSum_ready(dss_0_23_io_pSum_ready),
    .io_pSum_valid(dss_0_23_io_pSum_valid),
    .io_pSum_bits(dss_0_23_io_pSum_bits)
  );
  Node_25 NoC_1_0 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_0_clock),
    .reset(NoC_1_0_reset),
    .io_dataPackageIn_ready(NoC_1_0_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_0_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_0_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_0_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_row(NoC_1_0_io_dataPackageIn_bits_positon_row),
    .io_dataPackageIn_bits_positon_col(NoC_1_0_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_0_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_0_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_0_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_0_io_dataPackageOut_bits_dataType),
    .io_dataPackageOut_bits_positon_col(NoC_1_0_io_dataPackageOut_bits_positon_col)
  );
  Node_26 NoC_1_1 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_1_clock),
    .reset(NoC_1_1_reset),
    .io_dataPackageIn_ready(NoC_1_1_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_1_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_1_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_1_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_1_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_1_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_1_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_1_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_1_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_0 ( // @[PEArray.scala 36:24]
    .clock(pes_1_0_clock),
    .reset(pes_1_0_reset),
    .io_stateSW(pes_1_0_io_stateSW),
    .io_peconfig_ready(pes_1_0_io_peconfig_ready),
    .io_peconfig_valid(pes_1_0_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_0_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_0_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_0_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_0_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_0_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_0_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_0_io_filter_ready),
    .io_filter_valid(pes_1_0_io_filter_valid),
    .io_filter_bits(pes_1_0_io_filter_bits),
    .io_ifmap_ready(pes_1_0_io_ifmap_ready),
    .io_ifmap_valid(pes_1_0_io_ifmap_valid),
    .io_ifmap_bits(pes_1_0_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_0_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_0_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_0_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_0_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_0_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_0_io_pSumOut_bits),
    .io_stateOut(pes_1_0_io_stateOut)
  );
  dataSwitch dss_1_0 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_0_io_dataIn_ready),
    .io_dataIn_valid(dss_1_0_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_0_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_0_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_0_io_filter_ready),
    .io_filter_valid(dss_1_0_io_filter_valid),
    .io_filter_bits(dss_1_0_io_filter_bits),
    .io_ifmap_ready(dss_1_0_io_ifmap_ready),
    .io_ifmap_valid(dss_1_0_io_ifmap_valid),
    .io_ifmap_bits(dss_1_0_io_ifmap_bits),
    .io_pSum_ready(dss_1_0_io_pSum_ready),
    .io_pSum_valid(dss_1_0_io_pSum_valid),
    .io_pSum_bits(dss_1_0_io_pSum_bits)
  );
  Node_27 NoC_1_2 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_2_clock),
    .reset(NoC_1_2_reset),
    .io_dataPackageIn_ready(NoC_1_2_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_2_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_2_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_2_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_2_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_2_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_2_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_2_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_2_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_1 ( // @[PEArray.scala 36:24]
    .clock(pes_1_1_clock),
    .reset(pes_1_1_reset),
    .io_stateSW(pes_1_1_io_stateSW),
    .io_peconfig_ready(pes_1_1_io_peconfig_ready),
    .io_peconfig_valid(pes_1_1_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_1_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_1_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_1_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_1_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_1_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_1_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_1_io_filter_ready),
    .io_filter_valid(pes_1_1_io_filter_valid),
    .io_filter_bits(pes_1_1_io_filter_bits),
    .io_ifmap_ready(pes_1_1_io_ifmap_ready),
    .io_ifmap_valid(pes_1_1_io_ifmap_valid),
    .io_ifmap_bits(pes_1_1_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_1_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_1_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_1_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_1_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_1_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_1_io_pSumOut_bits),
    .io_stateOut(pes_1_1_io_stateOut)
  );
  dataSwitch dss_1_1 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_1_io_dataIn_ready),
    .io_dataIn_valid(dss_1_1_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_1_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_1_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_1_io_filter_ready),
    .io_filter_valid(dss_1_1_io_filter_valid),
    .io_filter_bits(dss_1_1_io_filter_bits),
    .io_ifmap_ready(dss_1_1_io_ifmap_ready),
    .io_ifmap_valid(dss_1_1_io_ifmap_valid),
    .io_ifmap_bits(dss_1_1_io_ifmap_bits),
    .io_pSum_ready(dss_1_1_io_pSum_ready),
    .io_pSum_valid(dss_1_1_io_pSum_valid),
    .io_pSum_bits(dss_1_1_io_pSum_bits)
  );
  Node_28 NoC_1_3 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_3_clock),
    .reset(NoC_1_3_reset),
    .io_dataPackageIn_ready(NoC_1_3_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_3_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_3_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_3_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_3_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_3_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_3_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_3_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_3_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_2 ( // @[PEArray.scala 36:24]
    .clock(pes_1_2_clock),
    .reset(pes_1_2_reset),
    .io_stateSW(pes_1_2_io_stateSW),
    .io_peconfig_ready(pes_1_2_io_peconfig_ready),
    .io_peconfig_valid(pes_1_2_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_2_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_2_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_2_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_2_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_2_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_2_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_2_io_filter_ready),
    .io_filter_valid(pes_1_2_io_filter_valid),
    .io_filter_bits(pes_1_2_io_filter_bits),
    .io_ifmap_ready(pes_1_2_io_ifmap_ready),
    .io_ifmap_valid(pes_1_2_io_ifmap_valid),
    .io_ifmap_bits(pes_1_2_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_2_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_2_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_2_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_2_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_2_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_2_io_pSumOut_bits),
    .io_stateOut(pes_1_2_io_stateOut)
  );
  dataSwitch dss_1_2 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_2_io_dataIn_ready),
    .io_dataIn_valid(dss_1_2_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_2_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_2_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_2_io_filter_ready),
    .io_filter_valid(dss_1_2_io_filter_valid),
    .io_filter_bits(dss_1_2_io_filter_bits),
    .io_ifmap_ready(dss_1_2_io_ifmap_ready),
    .io_ifmap_valid(dss_1_2_io_ifmap_valid),
    .io_ifmap_bits(dss_1_2_io_ifmap_bits),
    .io_pSum_ready(dss_1_2_io_pSum_ready),
    .io_pSum_valid(dss_1_2_io_pSum_valid),
    .io_pSum_bits(dss_1_2_io_pSum_bits)
  );
  Node_29 NoC_1_4 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_4_clock),
    .reset(NoC_1_4_reset),
    .io_dataPackageIn_ready(NoC_1_4_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_4_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_4_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_4_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_4_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_4_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_4_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_4_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_4_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_3 ( // @[PEArray.scala 36:24]
    .clock(pes_1_3_clock),
    .reset(pes_1_3_reset),
    .io_stateSW(pes_1_3_io_stateSW),
    .io_peconfig_ready(pes_1_3_io_peconfig_ready),
    .io_peconfig_valid(pes_1_3_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_3_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_3_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_3_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_3_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_3_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_3_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_3_io_filter_ready),
    .io_filter_valid(pes_1_3_io_filter_valid),
    .io_filter_bits(pes_1_3_io_filter_bits),
    .io_ifmap_ready(pes_1_3_io_ifmap_ready),
    .io_ifmap_valid(pes_1_3_io_ifmap_valid),
    .io_ifmap_bits(pes_1_3_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_3_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_3_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_3_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_3_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_3_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_3_io_pSumOut_bits),
    .io_stateOut(pes_1_3_io_stateOut)
  );
  dataSwitch dss_1_3 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_3_io_dataIn_ready),
    .io_dataIn_valid(dss_1_3_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_3_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_3_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_3_io_filter_ready),
    .io_filter_valid(dss_1_3_io_filter_valid),
    .io_filter_bits(dss_1_3_io_filter_bits),
    .io_ifmap_ready(dss_1_3_io_ifmap_ready),
    .io_ifmap_valid(dss_1_3_io_ifmap_valid),
    .io_ifmap_bits(dss_1_3_io_ifmap_bits),
    .io_pSum_ready(dss_1_3_io_pSum_ready),
    .io_pSum_valid(dss_1_3_io_pSum_valid),
    .io_pSum_bits(dss_1_3_io_pSum_bits)
  );
  Node_30 NoC_1_5 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_5_clock),
    .reset(NoC_1_5_reset),
    .io_dataPackageIn_ready(NoC_1_5_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_5_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_5_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_5_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_5_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_5_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_5_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_5_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_5_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_4 ( // @[PEArray.scala 36:24]
    .clock(pes_1_4_clock),
    .reset(pes_1_4_reset),
    .io_stateSW(pes_1_4_io_stateSW),
    .io_peconfig_ready(pes_1_4_io_peconfig_ready),
    .io_peconfig_valid(pes_1_4_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_4_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_4_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_4_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_4_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_4_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_4_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_4_io_filter_ready),
    .io_filter_valid(pes_1_4_io_filter_valid),
    .io_filter_bits(pes_1_4_io_filter_bits),
    .io_ifmap_ready(pes_1_4_io_ifmap_ready),
    .io_ifmap_valid(pes_1_4_io_ifmap_valid),
    .io_ifmap_bits(pes_1_4_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_4_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_4_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_4_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_4_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_4_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_4_io_pSumOut_bits),
    .io_stateOut(pes_1_4_io_stateOut)
  );
  dataSwitch dss_1_4 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_4_io_dataIn_ready),
    .io_dataIn_valid(dss_1_4_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_4_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_4_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_4_io_filter_ready),
    .io_filter_valid(dss_1_4_io_filter_valid),
    .io_filter_bits(dss_1_4_io_filter_bits),
    .io_ifmap_ready(dss_1_4_io_ifmap_ready),
    .io_ifmap_valid(dss_1_4_io_ifmap_valid),
    .io_ifmap_bits(dss_1_4_io_ifmap_bits),
    .io_pSum_ready(dss_1_4_io_pSum_ready),
    .io_pSum_valid(dss_1_4_io_pSum_valid),
    .io_pSum_bits(dss_1_4_io_pSum_bits)
  );
  Node_31 NoC_1_6 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_6_clock),
    .reset(NoC_1_6_reset),
    .io_dataPackageIn_ready(NoC_1_6_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_6_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_6_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_6_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_6_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_6_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_6_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_6_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_6_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_5 ( // @[PEArray.scala 36:24]
    .clock(pes_1_5_clock),
    .reset(pes_1_5_reset),
    .io_stateSW(pes_1_5_io_stateSW),
    .io_peconfig_ready(pes_1_5_io_peconfig_ready),
    .io_peconfig_valid(pes_1_5_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_5_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_5_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_5_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_5_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_5_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_5_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_5_io_filter_ready),
    .io_filter_valid(pes_1_5_io_filter_valid),
    .io_filter_bits(pes_1_5_io_filter_bits),
    .io_ifmap_ready(pes_1_5_io_ifmap_ready),
    .io_ifmap_valid(pes_1_5_io_ifmap_valid),
    .io_ifmap_bits(pes_1_5_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_5_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_5_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_5_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_5_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_5_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_5_io_pSumOut_bits),
    .io_stateOut(pes_1_5_io_stateOut)
  );
  dataSwitch dss_1_5 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_5_io_dataIn_ready),
    .io_dataIn_valid(dss_1_5_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_5_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_5_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_5_io_filter_ready),
    .io_filter_valid(dss_1_5_io_filter_valid),
    .io_filter_bits(dss_1_5_io_filter_bits),
    .io_ifmap_ready(dss_1_5_io_ifmap_ready),
    .io_ifmap_valid(dss_1_5_io_ifmap_valid),
    .io_ifmap_bits(dss_1_5_io_ifmap_bits),
    .io_pSum_ready(dss_1_5_io_pSum_ready),
    .io_pSum_valid(dss_1_5_io_pSum_valid),
    .io_pSum_bits(dss_1_5_io_pSum_bits)
  );
  Node_32 NoC_1_7 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_7_clock),
    .reset(NoC_1_7_reset),
    .io_dataPackageIn_ready(NoC_1_7_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_7_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_7_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_7_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_7_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_7_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_7_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_7_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_7_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_6 ( // @[PEArray.scala 36:24]
    .clock(pes_1_6_clock),
    .reset(pes_1_6_reset),
    .io_stateSW(pes_1_6_io_stateSW),
    .io_peconfig_ready(pes_1_6_io_peconfig_ready),
    .io_peconfig_valid(pes_1_6_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_6_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_6_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_6_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_6_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_6_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_6_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_6_io_filter_ready),
    .io_filter_valid(pes_1_6_io_filter_valid),
    .io_filter_bits(pes_1_6_io_filter_bits),
    .io_ifmap_ready(pes_1_6_io_ifmap_ready),
    .io_ifmap_valid(pes_1_6_io_ifmap_valid),
    .io_ifmap_bits(pes_1_6_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_6_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_6_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_6_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_6_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_6_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_6_io_pSumOut_bits),
    .io_stateOut(pes_1_6_io_stateOut)
  );
  dataSwitch dss_1_6 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_6_io_dataIn_ready),
    .io_dataIn_valid(dss_1_6_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_6_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_6_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_6_io_filter_ready),
    .io_filter_valid(dss_1_6_io_filter_valid),
    .io_filter_bits(dss_1_6_io_filter_bits),
    .io_ifmap_ready(dss_1_6_io_ifmap_ready),
    .io_ifmap_valid(dss_1_6_io_ifmap_valid),
    .io_ifmap_bits(dss_1_6_io_ifmap_bits),
    .io_pSum_ready(dss_1_6_io_pSum_ready),
    .io_pSum_valid(dss_1_6_io_pSum_valid),
    .io_pSum_bits(dss_1_6_io_pSum_bits)
  );
  Node_33 NoC_1_8 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_8_clock),
    .reset(NoC_1_8_reset),
    .io_dataPackageIn_ready(NoC_1_8_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_8_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_8_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_8_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_8_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_8_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_8_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_8_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_8_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_7 ( // @[PEArray.scala 36:24]
    .clock(pes_1_7_clock),
    .reset(pes_1_7_reset),
    .io_stateSW(pes_1_7_io_stateSW),
    .io_peconfig_ready(pes_1_7_io_peconfig_ready),
    .io_peconfig_valid(pes_1_7_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_7_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_7_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_7_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_7_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_7_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_7_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_7_io_filter_ready),
    .io_filter_valid(pes_1_7_io_filter_valid),
    .io_filter_bits(pes_1_7_io_filter_bits),
    .io_ifmap_ready(pes_1_7_io_ifmap_ready),
    .io_ifmap_valid(pes_1_7_io_ifmap_valid),
    .io_ifmap_bits(pes_1_7_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_7_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_7_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_7_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_7_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_7_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_7_io_pSumOut_bits),
    .io_stateOut(pes_1_7_io_stateOut)
  );
  dataSwitch dss_1_7 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_7_io_dataIn_ready),
    .io_dataIn_valid(dss_1_7_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_7_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_7_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_7_io_filter_ready),
    .io_filter_valid(dss_1_7_io_filter_valid),
    .io_filter_bits(dss_1_7_io_filter_bits),
    .io_ifmap_ready(dss_1_7_io_ifmap_ready),
    .io_ifmap_valid(dss_1_7_io_ifmap_valid),
    .io_ifmap_bits(dss_1_7_io_ifmap_bits),
    .io_pSum_ready(dss_1_7_io_pSum_ready),
    .io_pSum_valid(dss_1_7_io_pSum_valid),
    .io_pSum_bits(dss_1_7_io_pSum_bits)
  );
  Node_34 NoC_1_9 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_9_clock),
    .reset(NoC_1_9_reset),
    .io_dataPackageIn_ready(NoC_1_9_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_9_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_9_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_9_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_9_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_9_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_9_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_9_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_9_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_8 ( // @[PEArray.scala 36:24]
    .clock(pes_1_8_clock),
    .reset(pes_1_8_reset),
    .io_stateSW(pes_1_8_io_stateSW),
    .io_peconfig_ready(pes_1_8_io_peconfig_ready),
    .io_peconfig_valid(pes_1_8_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_8_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_8_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_8_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_8_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_8_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_8_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_8_io_filter_ready),
    .io_filter_valid(pes_1_8_io_filter_valid),
    .io_filter_bits(pes_1_8_io_filter_bits),
    .io_ifmap_ready(pes_1_8_io_ifmap_ready),
    .io_ifmap_valid(pes_1_8_io_ifmap_valid),
    .io_ifmap_bits(pes_1_8_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_8_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_8_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_8_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_8_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_8_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_8_io_pSumOut_bits),
    .io_stateOut(pes_1_8_io_stateOut)
  );
  dataSwitch dss_1_8 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_8_io_dataIn_ready),
    .io_dataIn_valid(dss_1_8_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_8_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_8_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_8_io_filter_ready),
    .io_filter_valid(dss_1_8_io_filter_valid),
    .io_filter_bits(dss_1_8_io_filter_bits),
    .io_ifmap_ready(dss_1_8_io_ifmap_ready),
    .io_ifmap_valid(dss_1_8_io_ifmap_valid),
    .io_ifmap_bits(dss_1_8_io_ifmap_bits),
    .io_pSum_ready(dss_1_8_io_pSum_ready),
    .io_pSum_valid(dss_1_8_io_pSum_valid),
    .io_pSum_bits(dss_1_8_io_pSum_bits)
  );
  Node_35 NoC_1_10 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_10_clock),
    .reset(NoC_1_10_reset),
    .io_dataPackageIn_ready(NoC_1_10_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_10_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_10_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_10_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_10_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_10_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_10_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_10_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_10_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_9 ( // @[PEArray.scala 36:24]
    .clock(pes_1_9_clock),
    .reset(pes_1_9_reset),
    .io_stateSW(pes_1_9_io_stateSW),
    .io_peconfig_ready(pes_1_9_io_peconfig_ready),
    .io_peconfig_valid(pes_1_9_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_9_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_9_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_9_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_9_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_9_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_9_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_9_io_filter_ready),
    .io_filter_valid(pes_1_9_io_filter_valid),
    .io_filter_bits(pes_1_9_io_filter_bits),
    .io_ifmap_ready(pes_1_9_io_ifmap_ready),
    .io_ifmap_valid(pes_1_9_io_ifmap_valid),
    .io_ifmap_bits(pes_1_9_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_9_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_9_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_9_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_9_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_9_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_9_io_pSumOut_bits),
    .io_stateOut(pes_1_9_io_stateOut)
  );
  dataSwitch dss_1_9 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_9_io_dataIn_ready),
    .io_dataIn_valid(dss_1_9_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_9_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_9_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_9_io_filter_ready),
    .io_filter_valid(dss_1_9_io_filter_valid),
    .io_filter_bits(dss_1_9_io_filter_bits),
    .io_ifmap_ready(dss_1_9_io_ifmap_ready),
    .io_ifmap_valid(dss_1_9_io_ifmap_valid),
    .io_ifmap_bits(dss_1_9_io_ifmap_bits),
    .io_pSum_ready(dss_1_9_io_pSum_ready),
    .io_pSum_valid(dss_1_9_io_pSum_valid),
    .io_pSum_bits(dss_1_9_io_pSum_bits)
  );
  Node_36 NoC_1_11 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_11_clock),
    .reset(NoC_1_11_reset),
    .io_dataPackageIn_ready(NoC_1_11_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_11_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_11_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_11_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_11_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_11_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_11_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_11_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_11_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_10 ( // @[PEArray.scala 36:24]
    .clock(pes_1_10_clock),
    .reset(pes_1_10_reset),
    .io_stateSW(pes_1_10_io_stateSW),
    .io_peconfig_ready(pes_1_10_io_peconfig_ready),
    .io_peconfig_valid(pes_1_10_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_10_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_10_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_10_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_10_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_10_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_10_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_10_io_filter_ready),
    .io_filter_valid(pes_1_10_io_filter_valid),
    .io_filter_bits(pes_1_10_io_filter_bits),
    .io_ifmap_ready(pes_1_10_io_ifmap_ready),
    .io_ifmap_valid(pes_1_10_io_ifmap_valid),
    .io_ifmap_bits(pes_1_10_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_10_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_10_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_10_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_10_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_10_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_10_io_pSumOut_bits),
    .io_stateOut(pes_1_10_io_stateOut)
  );
  dataSwitch dss_1_10 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_10_io_dataIn_ready),
    .io_dataIn_valid(dss_1_10_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_10_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_10_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_10_io_filter_ready),
    .io_filter_valid(dss_1_10_io_filter_valid),
    .io_filter_bits(dss_1_10_io_filter_bits),
    .io_ifmap_ready(dss_1_10_io_ifmap_ready),
    .io_ifmap_valid(dss_1_10_io_ifmap_valid),
    .io_ifmap_bits(dss_1_10_io_ifmap_bits),
    .io_pSum_ready(dss_1_10_io_pSum_ready),
    .io_pSum_valid(dss_1_10_io_pSum_valid),
    .io_pSum_bits(dss_1_10_io_pSum_bits)
  );
  Node_37 NoC_1_12 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_12_clock),
    .reset(NoC_1_12_reset),
    .io_dataPackageIn_ready(NoC_1_12_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_12_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_12_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_12_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_12_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_12_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_12_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_12_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_12_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_11 ( // @[PEArray.scala 36:24]
    .clock(pes_1_11_clock),
    .reset(pes_1_11_reset),
    .io_stateSW(pes_1_11_io_stateSW),
    .io_peconfig_ready(pes_1_11_io_peconfig_ready),
    .io_peconfig_valid(pes_1_11_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_11_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_11_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_11_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_11_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_11_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_11_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_11_io_filter_ready),
    .io_filter_valid(pes_1_11_io_filter_valid),
    .io_filter_bits(pes_1_11_io_filter_bits),
    .io_ifmap_ready(pes_1_11_io_ifmap_ready),
    .io_ifmap_valid(pes_1_11_io_ifmap_valid),
    .io_ifmap_bits(pes_1_11_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_11_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_11_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_11_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_11_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_11_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_11_io_pSumOut_bits),
    .io_stateOut(pes_1_11_io_stateOut)
  );
  dataSwitch dss_1_11 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_11_io_dataIn_ready),
    .io_dataIn_valid(dss_1_11_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_11_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_11_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_11_io_filter_ready),
    .io_filter_valid(dss_1_11_io_filter_valid),
    .io_filter_bits(dss_1_11_io_filter_bits),
    .io_ifmap_ready(dss_1_11_io_ifmap_ready),
    .io_ifmap_valid(dss_1_11_io_ifmap_valid),
    .io_ifmap_bits(dss_1_11_io_ifmap_bits),
    .io_pSum_ready(dss_1_11_io_pSum_ready),
    .io_pSum_valid(dss_1_11_io_pSum_valid),
    .io_pSum_bits(dss_1_11_io_pSum_bits)
  );
  Node_38 NoC_1_13 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_13_clock),
    .reset(NoC_1_13_reset),
    .io_dataPackageIn_ready(NoC_1_13_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_13_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_13_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_13_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_13_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_13_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_13_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_13_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_13_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_12 ( // @[PEArray.scala 36:24]
    .clock(pes_1_12_clock),
    .reset(pes_1_12_reset),
    .io_stateSW(pes_1_12_io_stateSW),
    .io_peconfig_ready(pes_1_12_io_peconfig_ready),
    .io_peconfig_valid(pes_1_12_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_12_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_12_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_12_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_12_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_12_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_12_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_12_io_filter_ready),
    .io_filter_valid(pes_1_12_io_filter_valid),
    .io_filter_bits(pes_1_12_io_filter_bits),
    .io_ifmap_ready(pes_1_12_io_ifmap_ready),
    .io_ifmap_valid(pes_1_12_io_ifmap_valid),
    .io_ifmap_bits(pes_1_12_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_12_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_12_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_12_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_12_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_12_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_12_io_pSumOut_bits),
    .io_stateOut(pes_1_12_io_stateOut)
  );
  dataSwitch dss_1_12 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_12_io_dataIn_ready),
    .io_dataIn_valid(dss_1_12_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_12_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_12_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_12_io_filter_ready),
    .io_filter_valid(dss_1_12_io_filter_valid),
    .io_filter_bits(dss_1_12_io_filter_bits),
    .io_ifmap_ready(dss_1_12_io_ifmap_ready),
    .io_ifmap_valid(dss_1_12_io_ifmap_valid),
    .io_ifmap_bits(dss_1_12_io_ifmap_bits),
    .io_pSum_ready(dss_1_12_io_pSum_ready),
    .io_pSum_valid(dss_1_12_io_pSum_valid),
    .io_pSum_bits(dss_1_12_io_pSum_bits)
  );
  Node_39 NoC_1_14 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_14_clock),
    .reset(NoC_1_14_reset),
    .io_dataPackageIn_ready(NoC_1_14_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_14_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_14_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_14_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_14_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_14_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_14_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_14_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_14_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_13 ( // @[PEArray.scala 36:24]
    .clock(pes_1_13_clock),
    .reset(pes_1_13_reset),
    .io_stateSW(pes_1_13_io_stateSW),
    .io_peconfig_ready(pes_1_13_io_peconfig_ready),
    .io_peconfig_valid(pes_1_13_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_13_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_13_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_13_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_13_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_13_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_13_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_13_io_filter_ready),
    .io_filter_valid(pes_1_13_io_filter_valid),
    .io_filter_bits(pes_1_13_io_filter_bits),
    .io_ifmap_ready(pes_1_13_io_ifmap_ready),
    .io_ifmap_valid(pes_1_13_io_ifmap_valid),
    .io_ifmap_bits(pes_1_13_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_13_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_13_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_13_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_13_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_13_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_13_io_pSumOut_bits),
    .io_stateOut(pes_1_13_io_stateOut)
  );
  dataSwitch dss_1_13 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_13_io_dataIn_ready),
    .io_dataIn_valid(dss_1_13_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_13_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_13_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_13_io_filter_ready),
    .io_filter_valid(dss_1_13_io_filter_valid),
    .io_filter_bits(dss_1_13_io_filter_bits),
    .io_ifmap_ready(dss_1_13_io_ifmap_ready),
    .io_ifmap_valid(dss_1_13_io_ifmap_valid),
    .io_ifmap_bits(dss_1_13_io_ifmap_bits),
    .io_pSum_ready(dss_1_13_io_pSum_ready),
    .io_pSum_valid(dss_1_13_io_pSum_valid),
    .io_pSum_bits(dss_1_13_io_pSum_bits)
  );
  Node_40 NoC_1_15 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_15_clock),
    .reset(NoC_1_15_reset),
    .io_dataPackageIn_ready(NoC_1_15_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_15_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_15_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_15_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_15_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_15_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_15_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_15_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_15_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_14 ( // @[PEArray.scala 36:24]
    .clock(pes_1_14_clock),
    .reset(pes_1_14_reset),
    .io_stateSW(pes_1_14_io_stateSW),
    .io_peconfig_ready(pes_1_14_io_peconfig_ready),
    .io_peconfig_valid(pes_1_14_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_14_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_14_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_14_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_14_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_14_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_14_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_14_io_filter_ready),
    .io_filter_valid(pes_1_14_io_filter_valid),
    .io_filter_bits(pes_1_14_io_filter_bits),
    .io_ifmap_ready(pes_1_14_io_ifmap_ready),
    .io_ifmap_valid(pes_1_14_io_ifmap_valid),
    .io_ifmap_bits(pes_1_14_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_14_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_14_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_14_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_14_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_14_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_14_io_pSumOut_bits),
    .io_stateOut(pes_1_14_io_stateOut)
  );
  dataSwitch dss_1_14 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_14_io_dataIn_ready),
    .io_dataIn_valid(dss_1_14_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_14_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_14_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_14_io_filter_ready),
    .io_filter_valid(dss_1_14_io_filter_valid),
    .io_filter_bits(dss_1_14_io_filter_bits),
    .io_ifmap_ready(dss_1_14_io_ifmap_ready),
    .io_ifmap_valid(dss_1_14_io_ifmap_valid),
    .io_ifmap_bits(dss_1_14_io_ifmap_bits),
    .io_pSum_ready(dss_1_14_io_pSum_ready),
    .io_pSum_valid(dss_1_14_io_pSum_valid),
    .io_pSum_bits(dss_1_14_io_pSum_bits)
  );
  Node_41 NoC_1_16 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_16_clock),
    .reset(NoC_1_16_reset),
    .io_dataPackageIn_ready(NoC_1_16_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_16_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_16_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_16_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_16_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_16_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_16_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_16_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_16_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_15 ( // @[PEArray.scala 36:24]
    .clock(pes_1_15_clock),
    .reset(pes_1_15_reset),
    .io_stateSW(pes_1_15_io_stateSW),
    .io_peconfig_ready(pes_1_15_io_peconfig_ready),
    .io_peconfig_valid(pes_1_15_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_15_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_15_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_15_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_15_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_15_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_15_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_15_io_filter_ready),
    .io_filter_valid(pes_1_15_io_filter_valid),
    .io_filter_bits(pes_1_15_io_filter_bits),
    .io_ifmap_ready(pes_1_15_io_ifmap_ready),
    .io_ifmap_valid(pes_1_15_io_ifmap_valid),
    .io_ifmap_bits(pes_1_15_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_15_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_15_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_15_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_15_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_15_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_15_io_pSumOut_bits),
    .io_stateOut(pes_1_15_io_stateOut)
  );
  dataSwitch dss_1_15 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_15_io_dataIn_ready),
    .io_dataIn_valid(dss_1_15_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_15_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_15_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_15_io_filter_ready),
    .io_filter_valid(dss_1_15_io_filter_valid),
    .io_filter_bits(dss_1_15_io_filter_bits),
    .io_ifmap_ready(dss_1_15_io_ifmap_ready),
    .io_ifmap_valid(dss_1_15_io_ifmap_valid),
    .io_ifmap_bits(dss_1_15_io_ifmap_bits),
    .io_pSum_ready(dss_1_15_io_pSum_ready),
    .io_pSum_valid(dss_1_15_io_pSum_valid),
    .io_pSum_bits(dss_1_15_io_pSum_bits)
  );
  Node_42 NoC_1_17 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_17_clock),
    .reset(NoC_1_17_reset),
    .io_dataPackageIn_ready(NoC_1_17_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_17_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_17_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_17_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_17_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_17_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_17_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_17_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_17_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_16 ( // @[PEArray.scala 36:24]
    .clock(pes_1_16_clock),
    .reset(pes_1_16_reset),
    .io_stateSW(pes_1_16_io_stateSW),
    .io_peconfig_ready(pes_1_16_io_peconfig_ready),
    .io_peconfig_valid(pes_1_16_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_16_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_16_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_16_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_16_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_16_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_16_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_16_io_filter_ready),
    .io_filter_valid(pes_1_16_io_filter_valid),
    .io_filter_bits(pes_1_16_io_filter_bits),
    .io_ifmap_ready(pes_1_16_io_ifmap_ready),
    .io_ifmap_valid(pes_1_16_io_ifmap_valid),
    .io_ifmap_bits(pes_1_16_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_16_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_16_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_16_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_16_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_16_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_16_io_pSumOut_bits),
    .io_stateOut(pes_1_16_io_stateOut)
  );
  dataSwitch dss_1_16 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_16_io_dataIn_ready),
    .io_dataIn_valid(dss_1_16_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_16_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_16_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_16_io_filter_ready),
    .io_filter_valid(dss_1_16_io_filter_valid),
    .io_filter_bits(dss_1_16_io_filter_bits),
    .io_ifmap_ready(dss_1_16_io_ifmap_ready),
    .io_ifmap_valid(dss_1_16_io_ifmap_valid),
    .io_ifmap_bits(dss_1_16_io_ifmap_bits),
    .io_pSum_ready(dss_1_16_io_pSum_ready),
    .io_pSum_valid(dss_1_16_io_pSum_valid),
    .io_pSum_bits(dss_1_16_io_pSum_bits)
  );
  Node_43 NoC_1_18 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_18_clock),
    .reset(NoC_1_18_reset),
    .io_dataPackageIn_ready(NoC_1_18_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_18_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_18_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_18_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_18_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_18_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_18_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_18_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_18_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_17 ( // @[PEArray.scala 36:24]
    .clock(pes_1_17_clock),
    .reset(pes_1_17_reset),
    .io_stateSW(pes_1_17_io_stateSW),
    .io_peconfig_ready(pes_1_17_io_peconfig_ready),
    .io_peconfig_valid(pes_1_17_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_17_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_17_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_17_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_17_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_17_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_17_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_17_io_filter_ready),
    .io_filter_valid(pes_1_17_io_filter_valid),
    .io_filter_bits(pes_1_17_io_filter_bits),
    .io_ifmap_ready(pes_1_17_io_ifmap_ready),
    .io_ifmap_valid(pes_1_17_io_ifmap_valid),
    .io_ifmap_bits(pes_1_17_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_17_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_17_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_17_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_17_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_17_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_17_io_pSumOut_bits),
    .io_stateOut(pes_1_17_io_stateOut)
  );
  dataSwitch dss_1_17 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_17_io_dataIn_ready),
    .io_dataIn_valid(dss_1_17_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_17_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_17_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_17_io_filter_ready),
    .io_filter_valid(dss_1_17_io_filter_valid),
    .io_filter_bits(dss_1_17_io_filter_bits),
    .io_ifmap_ready(dss_1_17_io_ifmap_ready),
    .io_ifmap_valid(dss_1_17_io_ifmap_valid),
    .io_ifmap_bits(dss_1_17_io_ifmap_bits),
    .io_pSum_ready(dss_1_17_io_pSum_ready),
    .io_pSum_valid(dss_1_17_io_pSum_valid),
    .io_pSum_bits(dss_1_17_io_pSum_bits)
  );
  Node_44 NoC_1_19 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_19_clock),
    .reset(NoC_1_19_reset),
    .io_dataPackageIn_ready(NoC_1_19_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_19_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_19_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_19_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_19_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_19_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_19_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_19_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_19_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_18 ( // @[PEArray.scala 36:24]
    .clock(pes_1_18_clock),
    .reset(pes_1_18_reset),
    .io_stateSW(pes_1_18_io_stateSW),
    .io_peconfig_ready(pes_1_18_io_peconfig_ready),
    .io_peconfig_valid(pes_1_18_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_18_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_18_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_18_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_18_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_18_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_18_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_18_io_filter_ready),
    .io_filter_valid(pes_1_18_io_filter_valid),
    .io_filter_bits(pes_1_18_io_filter_bits),
    .io_ifmap_ready(pes_1_18_io_ifmap_ready),
    .io_ifmap_valid(pes_1_18_io_ifmap_valid),
    .io_ifmap_bits(pes_1_18_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_18_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_18_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_18_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_18_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_18_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_18_io_pSumOut_bits),
    .io_stateOut(pes_1_18_io_stateOut)
  );
  dataSwitch dss_1_18 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_18_io_dataIn_ready),
    .io_dataIn_valid(dss_1_18_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_18_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_18_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_18_io_filter_ready),
    .io_filter_valid(dss_1_18_io_filter_valid),
    .io_filter_bits(dss_1_18_io_filter_bits),
    .io_ifmap_ready(dss_1_18_io_ifmap_ready),
    .io_ifmap_valid(dss_1_18_io_ifmap_valid),
    .io_ifmap_bits(dss_1_18_io_ifmap_bits),
    .io_pSum_ready(dss_1_18_io_pSum_ready),
    .io_pSum_valid(dss_1_18_io_pSum_valid),
    .io_pSum_bits(dss_1_18_io_pSum_bits)
  );
  Node_45 NoC_1_20 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_20_clock),
    .reset(NoC_1_20_reset),
    .io_dataPackageIn_ready(NoC_1_20_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_20_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_20_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_20_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_20_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_20_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_20_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_20_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_20_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_19 ( // @[PEArray.scala 36:24]
    .clock(pes_1_19_clock),
    .reset(pes_1_19_reset),
    .io_stateSW(pes_1_19_io_stateSW),
    .io_peconfig_ready(pes_1_19_io_peconfig_ready),
    .io_peconfig_valid(pes_1_19_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_19_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_19_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_19_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_19_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_19_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_19_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_19_io_filter_ready),
    .io_filter_valid(pes_1_19_io_filter_valid),
    .io_filter_bits(pes_1_19_io_filter_bits),
    .io_ifmap_ready(pes_1_19_io_ifmap_ready),
    .io_ifmap_valid(pes_1_19_io_ifmap_valid),
    .io_ifmap_bits(pes_1_19_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_19_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_19_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_19_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_19_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_19_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_19_io_pSumOut_bits),
    .io_stateOut(pes_1_19_io_stateOut)
  );
  dataSwitch dss_1_19 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_19_io_dataIn_ready),
    .io_dataIn_valid(dss_1_19_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_19_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_19_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_19_io_filter_ready),
    .io_filter_valid(dss_1_19_io_filter_valid),
    .io_filter_bits(dss_1_19_io_filter_bits),
    .io_ifmap_ready(dss_1_19_io_ifmap_ready),
    .io_ifmap_valid(dss_1_19_io_ifmap_valid),
    .io_ifmap_bits(dss_1_19_io_ifmap_bits),
    .io_pSum_ready(dss_1_19_io_pSum_ready),
    .io_pSum_valid(dss_1_19_io_pSum_valid),
    .io_pSum_bits(dss_1_19_io_pSum_bits)
  );
  Node_46 NoC_1_21 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_21_clock),
    .reset(NoC_1_21_reset),
    .io_dataPackageIn_ready(NoC_1_21_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_21_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_21_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_21_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_21_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_21_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_21_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_21_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_21_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_20 ( // @[PEArray.scala 36:24]
    .clock(pes_1_20_clock),
    .reset(pes_1_20_reset),
    .io_stateSW(pes_1_20_io_stateSW),
    .io_peconfig_ready(pes_1_20_io_peconfig_ready),
    .io_peconfig_valid(pes_1_20_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_20_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_20_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_20_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_20_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_20_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_20_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_20_io_filter_ready),
    .io_filter_valid(pes_1_20_io_filter_valid),
    .io_filter_bits(pes_1_20_io_filter_bits),
    .io_ifmap_ready(pes_1_20_io_ifmap_ready),
    .io_ifmap_valid(pes_1_20_io_ifmap_valid),
    .io_ifmap_bits(pes_1_20_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_20_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_20_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_20_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_20_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_20_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_20_io_pSumOut_bits),
    .io_stateOut(pes_1_20_io_stateOut)
  );
  dataSwitch dss_1_20 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_20_io_dataIn_ready),
    .io_dataIn_valid(dss_1_20_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_20_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_20_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_20_io_filter_ready),
    .io_filter_valid(dss_1_20_io_filter_valid),
    .io_filter_bits(dss_1_20_io_filter_bits),
    .io_ifmap_ready(dss_1_20_io_ifmap_ready),
    .io_ifmap_valid(dss_1_20_io_ifmap_valid),
    .io_ifmap_bits(dss_1_20_io_ifmap_bits),
    .io_pSum_ready(dss_1_20_io_pSum_ready),
    .io_pSum_valid(dss_1_20_io_pSum_valid),
    .io_pSum_bits(dss_1_20_io_pSum_bits)
  );
  Node_47 NoC_1_22 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_22_clock),
    .reset(NoC_1_22_reset),
    .io_dataPackageIn_ready(NoC_1_22_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_22_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_22_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_22_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_22_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_22_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_22_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_22_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_22_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_21 ( // @[PEArray.scala 36:24]
    .clock(pes_1_21_clock),
    .reset(pes_1_21_reset),
    .io_stateSW(pes_1_21_io_stateSW),
    .io_peconfig_ready(pes_1_21_io_peconfig_ready),
    .io_peconfig_valid(pes_1_21_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_21_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_21_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_21_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_21_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_21_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_21_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_21_io_filter_ready),
    .io_filter_valid(pes_1_21_io_filter_valid),
    .io_filter_bits(pes_1_21_io_filter_bits),
    .io_ifmap_ready(pes_1_21_io_ifmap_ready),
    .io_ifmap_valid(pes_1_21_io_ifmap_valid),
    .io_ifmap_bits(pes_1_21_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_21_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_21_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_21_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_21_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_21_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_21_io_pSumOut_bits),
    .io_stateOut(pes_1_21_io_stateOut)
  );
  dataSwitch dss_1_21 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_21_io_dataIn_ready),
    .io_dataIn_valid(dss_1_21_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_21_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_21_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_21_io_filter_ready),
    .io_filter_valid(dss_1_21_io_filter_valid),
    .io_filter_bits(dss_1_21_io_filter_bits),
    .io_ifmap_ready(dss_1_21_io_ifmap_ready),
    .io_ifmap_valid(dss_1_21_io_ifmap_valid),
    .io_ifmap_bits(dss_1_21_io_ifmap_bits),
    .io_pSum_ready(dss_1_21_io_pSum_ready),
    .io_pSum_valid(dss_1_21_io_pSum_valid),
    .io_pSum_bits(dss_1_21_io_pSum_bits)
  );
  Node_48 NoC_1_23 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_23_clock),
    .reset(NoC_1_23_reset),
    .io_dataPackageIn_ready(NoC_1_23_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_23_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_23_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_23_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_23_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_23_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_23_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_23_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_23_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_22 ( // @[PEArray.scala 36:24]
    .clock(pes_1_22_clock),
    .reset(pes_1_22_reset),
    .io_stateSW(pes_1_22_io_stateSW),
    .io_peconfig_ready(pes_1_22_io_peconfig_ready),
    .io_peconfig_valid(pes_1_22_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_22_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_22_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_22_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_22_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_22_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_22_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_22_io_filter_ready),
    .io_filter_valid(pes_1_22_io_filter_valid),
    .io_filter_bits(pes_1_22_io_filter_bits),
    .io_ifmap_ready(pes_1_22_io_ifmap_ready),
    .io_ifmap_valid(pes_1_22_io_ifmap_valid),
    .io_ifmap_bits(pes_1_22_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_22_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_22_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_22_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_22_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_22_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_22_io_pSumOut_bits),
    .io_stateOut(pes_1_22_io_stateOut)
  );
  dataSwitch dss_1_22 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_22_io_dataIn_ready),
    .io_dataIn_valid(dss_1_22_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_22_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_22_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_22_io_filter_ready),
    .io_filter_valid(dss_1_22_io_filter_valid),
    .io_filter_bits(dss_1_22_io_filter_bits),
    .io_ifmap_ready(dss_1_22_io_ifmap_ready),
    .io_ifmap_valid(dss_1_22_io_ifmap_valid),
    .io_ifmap_bits(dss_1_22_io_ifmap_bits),
    .io_pSum_ready(dss_1_22_io_pSum_ready),
    .io_pSum_valid(dss_1_22_io_pSum_valid),
    .io_pSum_bits(dss_1_22_io_pSum_bits)
  );
  Node_49 NoC_1_24 ( // @[PEArray.scala 34:24]
    .clock(NoC_1_24_clock),
    .reset(NoC_1_24_reset),
    .io_dataPackageIn_ready(NoC_1_24_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_1_24_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_1_24_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_1_24_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_1_24_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_1_24_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_1_24_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_1_24_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_1_24_io_dataPackageOut_bits_dataType)
  );
  PETop pes_1_23 ( // @[PEArray.scala 36:24]
    .clock(pes_1_23_clock),
    .reset(pes_1_23_reset),
    .io_stateSW(pes_1_23_io_stateSW),
    .io_peconfig_ready(pes_1_23_io_peconfig_ready),
    .io_peconfig_valid(pes_1_23_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_1_23_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_1_23_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_1_23_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_1_23_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_1_23_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_1_23_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_1_23_io_filter_ready),
    .io_filter_valid(pes_1_23_io_filter_valid),
    .io_filter_bits(pes_1_23_io_filter_bits),
    .io_ifmap_ready(pes_1_23_io_ifmap_ready),
    .io_ifmap_valid(pes_1_23_io_ifmap_valid),
    .io_ifmap_bits(pes_1_23_io_ifmap_bits),
    .io_pSumIn_ready(pes_1_23_io_pSumIn_ready),
    .io_pSumIn_valid(pes_1_23_io_pSumIn_valid),
    .io_pSumIn_bits(pes_1_23_io_pSumIn_bits),
    .io_pSumOut_ready(pes_1_23_io_pSumOut_ready),
    .io_pSumOut_valid(pes_1_23_io_pSumOut_valid),
    .io_pSumOut_bits(pes_1_23_io_pSumOut_bits),
    .io_stateOut(pes_1_23_io_stateOut)
  );
  dataSwitch dss_1_23 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_1_23_io_dataIn_ready),
    .io_dataIn_valid(dss_1_23_io_dataIn_valid),
    .io_dataIn_bits_data(dss_1_23_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_1_23_io_dataIn_bits_dataType),
    .io_filter_ready(dss_1_23_io_filter_ready),
    .io_filter_valid(dss_1_23_io_filter_valid),
    .io_filter_bits(dss_1_23_io_filter_bits),
    .io_ifmap_ready(dss_1_23_io_ifmap_ready),
    .io_ifmap_valid(dss_1_23_io_ifmap_valid),
    .io_ifmap_bits(dss_1_23_io_ifmap_bits),
    .io_pSum_ready(dss_1_23_io_pSum_ready),
    .io_pSum_valid(dss_1_23_io_pSum_valid),
    .io_pSum_bits(dss_1_23_io_pSum_bits)
  );
  Node_50 NoC_2_0 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_0_clock),
    .reset(NoC_2_0_reset),
    .io_dataPackageIn_ready(NoC_2_0_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_0_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_0_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_0_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_row(NoC_2_0_io_dataPackageIn_bits_positon_row),
    .io_dataPackageIn_bits_positon_col(NoC_2_0_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_0_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_0_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_0_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_0_io_dataPackageOut_bits_dataType),
    .io_dataPackageOut_bits_positon_col(NoC_2_0_io_dataPackageOut_bits_positon_col)
  );
  Node_51 NoC_2_1 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_1_clock),
    .reset(NoC_2_1_reset),
    .io_dataPackageIn_ready(NoC_2_1_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_1_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_1_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_1_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_1_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_1_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_1_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_1_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_1_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_0 ( // @[PEArray.scala 36:24]
    .clock(pes_2_0_clock),
    .reset(pes_2_0_reset),
    .io_stateSW(pes_2_0_io_stateSW),
    .io_peconfig_ready(pes_2_0_io_peconfig_ready),
    .io_peconfig_valid(pes_2_0_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_0_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_0_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_0_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_0_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_0_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_0_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_0_io_filter_ready),
    .io_filter_valid(pes_2_0_io_filter_valid),
    .io_filter_bits(pes_2_0_io_filter_bits),
    .io_ifmap_ready(pes_2_0_io_ifmap_ready),
    .io_ifmap_valid(pes_2_0_io_ifmap_valid),
    .io_ifmap_bits(pes_2_0_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_0_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_0_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_0_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_0_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_0_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_0_io_pSumOut_bits),
    .io_stateOut(pes_2_0_io_stateOut)
  );
  dataSwitch dss_2_0 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_0_io_dataIn_ready),
    .io_dataIn_valid(dss_2_0_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_0_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_0_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_0_io_filter_ready),
    .io_filter_valid(dss_2_0_io_filter_valid),
    .io_filter_bits(dss_2_0_io_filter_bits),
    .io_ifmap_ready(dss_2_0_io_ifmap_ready),
    .io_ifmap_valid(dss_2_0_io_ifmap_valid),
    .io_ifmap_bits(dss_2_0_io_ifmap_bits),
    .io_pSum_ready(dss_2_0_io_pSum_ready),
    .io_pSum_valid(dss_2_0_io_pSum_valid),
    .io_pSum_bits(dss_2_0_io_pSum_bits)
  );
  Node_52 NoC_2_2 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_2_clock),
    .reset(NoC_2_2_reset),
    .io_dataPackageIn_ready(NoC_2_2_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_2_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_2_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_2_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_2_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_2_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_2_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_2_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_2_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_1 ( // @[PEArray.scala 36:24]
    .clock(pes_2_1_clock),
    .reset(pes_2_1_reset),
    .io_stateSW(pes_2_1_io_stateSW),
    .io_peconfig_ready(pes_2_1_io_peconfig_ready),
    .io_peconfig_valid(pes_2_1_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_1_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_1_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_1_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_1_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_1_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_1_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_1_io_filter_ready),
    .io_filter_valid(pes_2_1_io_filter_valid),
    .io_filter_bits(pes_2_1_io_filter_bits),
    .io_ifmap_ready(pes_2_1_io_ifmap_ready),
    .io_ifmap_valid(pes_2_1_io_ifmap_valid),
    .io_ifmap_bits(pes_2_1_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_1_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_1_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_1_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_1_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_1_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_1_io_pSumOut_bits),
    .io_stateOut(pes_2_1_io_stateOut)
  );
  dataSwitch dss_2_1 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_1_io_dataIn_ready),
    .io_dataIn_valid(dss_2_1_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_1_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_1_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_1_io_filter_ready),
    .io_filter_valid(dss_2_1_io_filter_valid),
    .io_filter_bits(dss_2_1_io_filter_bits),
    .io_ifmap_ready(dss_2_1_io_ifmap_ready),
    .io_ifmap_valid(dss_2_1_io_ifmap_valid),
    .io_ifmap_bits(dss_2_1_io_ifmap_bits),
    .io_pSum_ready(dss_2_1_io_pSum_ready),
    .io_pSum_valid(dss_2_1_io_pSum_valid),
    .io_pSum_bits(dss_2_1_io_pSum_bits)
  );
  Node_53 NoC_2_3 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_3_clock),
    .reset(NoC_2_3_reset),
    .io_dataPackageIn_ready(NoC_2_3_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_3_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_3_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_3_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_3_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_3_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_3_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_3_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_3_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_2 ( // @[PEArray.scala 36:24]
    .clock(pes_2_2_clock),
    .reset(pes_2_2_reset),
    .io_stateSW(pes_2_2_io_stateSW),
    .io_peconfig_ready(pes_2_2_io_peconfig_ready),
    .io_peconfig_valid(pes_2_2_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_2_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_2_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_2_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_2_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_2_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_2_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_2_io_filter_ready),
    .io_filter_valid(pes_2_2_io_filter_valid),
    .io_filter_bits(pes_2_2_io_filter_bits),
    .io_ifmap_ready(pes_2_2_io_ifmap_ready),
    .io_ifmap_valid(pes_2_2_io_ifmap_valid),
    .io_ifmap_bits(pes_2_2_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_2_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_2_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_2_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_2_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_2_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_2_io_pSumOut_bits),
    .io_stateOut(pes_2_2_io_stateOut)
  );
  dataSwitch dss_2_2 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_2_io_dataIn_ready),
    .io_dataIn_valid(dss_2_2_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_2_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_2_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_2_io_filter_ready),
    .io_filter_valid(dss_2_2_io_filter_valid),
    .io_filter_bits(dss_2_2_io_filter_bits),
    .io_ifmap_ready(dss_2_2_io_ifmap_ready),
    .io_ifmap_valid(dss_2_2_io_ifmap_valid),
    .io_ifmap_bits(dss_2_2_io_ifmap_bits),
    .io_pSum_ready(dss_2_2_io_pSum_ready),
    .io_pSum_valid(dss_2_2_io_pSum_valid),
    .io_pSum_bits(dss_2_2_io_pSum_bits)
  );
  Node_54 NoC_2_4 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_4_clock),
    .reset(NoC_2_4_reset),
    .io_dataPackageIn_ready(NoC_2_4_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_4_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_4_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_4_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_4_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_4_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_4_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_4_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_4_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_3 ( // @[PEArray.scala 36:24]
    .clock(pes_2_3_clock),
    .reset(pes_2_3_reset),
    .io_stateSW(pes_2_3_io_stateSW),
    .io_peconfig_ready(pes_2_3_io_peconfig_ready),
    .io_peconfig_valid(pes_2_3_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_3_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_3_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_3_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_3_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_3_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_3_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_3_io_filter_ready),
    .io_filter_valid(pes_2_3_io_filter_valid),
    .io_filter_bits(pes_2_3_io_filter_bits),
    .io_ifmap_ready(pes_2_3_io_ifmap_ready),
    .io_ifmap_valid(pes_2_3_io_ifmap_valid),
    .io_ifmap_bits(pes_2_3_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_3_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_3_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_3_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_3_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_3_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_3_io_pSumOut_bits),
    .io_stateOut(pes_2_3_io_stateOut)
  );
  dataSwitch dss_2_3 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_3_io_dataIn_ready),
    .io_dataIn_valid(dss_2_3_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_3_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_3_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_3_io_filter_ready),
    .io_filter_valid(dss_2_3_io_filter_valid),
    .io_filter_bits(dss_2_3_io_filter_bits),
    .io_ifmap_ready(dss_2_3_io_ifmap_ready),
    .io_ifmap_valid(dss_2_3_io_ifmap_valid),
    .io_ifmap_bits(dss_2_3_io_ifmap_bits),
    .io_pSum_ready(dss_2_3_io_pSum_ready),
    .io_pSum_valid(dss_2_3_io_pSum_valid),
    .io_pSum_bits(dss_2_3_io_pSum_bits)
  );
  Node_55 NoC_2_5 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_5_clock),
    .reset(NoC_2_5_reset),
    .io_dataPackageIn_ready(NoC_2_5_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_5_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_5_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_5_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_5_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_5_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_5_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_5_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_5_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_4 ( // @[PEArray.scala 36:24]
    .clock(pes_2_4_clock),
    .reset(pes_2_4_reset),
    .io_stateSW(pes_2_4_io_stateSW),
    .io_peconfig_ready(pes_2_4_io_peconfig_ready),
    .io_peconfig_valid(pes_2_4_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_4_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_4_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_4_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_4_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_4_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_4_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_4_io_filter_ready),
    .io_filter_valid(pes_2_4_io_filter_valid),
    .io_filter_bits(pes_2_4_io_filter_bits),
    .io_ifmap_ready(pes_2_4_io_ifmap_ready),
    .io_ifmap_valid(pes_2_4_io_ifmap_valid),
    .io_ifmap_bits(pes_2_4_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_4_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_4_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_4_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_4_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_4_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_4_io_pSumOut_bits),
    .io_stateOut(pes_2_4_io_stateOut)
  );
  dataSwitch dss_2_4 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_4_io_dataIn_ready),
    .io_dataIn_valid(dss_2_4_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_4_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_4_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_4_io_filter_ready),
    .io_filter_valid(dss_2_4_io_filter_valid),
    .io_filter_bits(dss_2_4_io_filter_bits),
    .io_ifmap_ready(dss_2_4_io_ifmap_ready),
    .io_ifmap_valid(dss_2_4_io_ifmap_valid),
    .io_ifmap_bits(dss_2_4_io_ifmap_bits),
    .io_pSum_ready(dss_2_4_io_pSum_ready),
    .io_pSum_valid(dss_2_4_io_pSum_valid),
    .io_pSum_bits(dss_2_4_io_pSum_bits)
  );
  Node_56 NoC_2_6 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_6_clock),
    .reset(NoC_2_6_reset),
    .io_dataPackageIn_ready(NoC_2_6_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_6_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_6_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_6_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_6_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_6_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_6_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_6_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_6_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_5 ( // @[PEArray.scala 36:24]
    .clock(pes_2_5_clock),
    .reset(pes_2_5_reset),
    .io_stateSW(pes_2_5_io_stateSW),
    .io_peconfig_ready(pes_2_5_io_peconfig_ready),
    .io_peconfig_valid(pes_2_5_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_5_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_5_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_5_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_5_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_5_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_5_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_5_io_filter_ready),
    .io_filter_valid(pes_2_5_io_filter_valid),
    .io_filter_bits(pes_2_5_io_filter_bits),
    .io_ifmap_ready(pes_2_5_io_ifmap_ready),
    .io_ifmap_valid(pes_2_5_io_ifmap_valid),
    .io_ifmap_bits(pes_2_5_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_5_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_5_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_5_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_5_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_5_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_5_io_pSumOut_bits),
    .io_stateOut(pes_2_5_io_stateOut)
  );
  dataSwitch dss_2_5 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_5_io_dataIn_ready),
    .io_dataIn_valid(dss_2_5_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_5_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_5_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_5_io_filter_ready),
    .io_filter_valid(dss_2_5_io_filter_valid),
    .io_filter_bits(dss_2_5_io_filter_bits),
    .io_ifmap_ready(dss_2_5_io_ifmap_ready),
    .io_ifmap_valid(dss_2_5_io_ifmap_valid),
    .io_ifmap_bits(dss_2_5_io_ifmap_bits),
    .io_pSum_ready(dss_2_5_io_pSum_ready),
    .io_pSum_valid(dss_2_5_io_pSum_valid),
    .io_pSum_bits(dss_2_5_io_pSum_bits)
  );
  Node_57 NoC_2_7 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_7_clock),
    .reset(NoC_2_7_reset),
    .io_dataPackageIn_ready(NoC_2_7_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_7_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_7_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_7_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_7_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_7_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_7_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_7_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_7_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_6 ( // @[PEArray.scala 36:24]
    .clock(pes_2_6_clock),
    .reset(pes_2_6_reset),
    .io_stateSW(pes_2_6_io_stateSW),
    .io_peconfig_ready(pes_2_6_io_peconfig_ready),
    .io_peconfig_valid(pes_2_6_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_6_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_6_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_6_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_6_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_6_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_6_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_6_io_filter_ready),
    .io_filter_valid(pes_2_6_io_filter_valid),
    .io_filter_bits(pes_2_6_io_filter_bits),
    .io_ifmap_ready(pes_2_6_io_ifmap_ready),
    .io_ifmap_valid(pes_2_6_io_ifmap_valid),
    .io_ifmap_bits(pes_2_6_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_6_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_6_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_6_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_6_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_6_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_6_io_pSumOut_bits),
    .io_stateOut(pes_2_6_io_stateOut)
  );
  dataSwitch dss_2_6 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_6_io_dataIn_ready),
    .io_dataIn_valid(dss_2_6_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_6_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_6_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_6_io_filter_ready),
    .io_filter_valid(dss_2_6_io_filter_valid),
    .io_filter_bits(dss_2_6_io_filter_bits),
    .io_ifmap_ready(dss_2_6_io_ifmap_ready),
    .io_ifmap_valid(dss_2_6_io_ifmap_valid),
    .io_ifmap_bits(dss_2_6_io_ifmap_bits),
    .io_pSum_ready(dss_2_6_io_pSum_ready),
    .io_pSum_valid(dss_2_6_io_pSum_valid),
    .io_pSum_bits(dss_2_6_io_pSum_bits)
  );
  Node_58 NoC_2_8 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_8_clock),
    .reset(NoC_2_8_reset),
    .io_dataPackageIn_ready(NoC_2_8_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_8_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_8_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_8_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_8_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_8_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_8_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_8_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_8_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_7 ( // @[PEArray.scala 36:24]
    .clock(pes_2_7_clock),
    .reset(pes_2_7_reset),
    .io_stateSW(pes_2_7_io_stateSW),
    .io_peconfig_ready(pes_2_7_io_peconfig_ready),
    .io_peconfig_valid(pes_2_7_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_7_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_7_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_7_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_7_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_7_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_7_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_7_io_filter_ready),
    .io_filter_valid(pes_2_7_io_filter_valid),
    .io_filter_bits(pes_2_7_io_filter_bits),
    .io_ifmap_ready(pes_2_7_io_ifmap_ready),
    .io_ifmap_valid(pes_2_7_io_ifmap_valid),
    .io_ifmap_bits(pes_2_7_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_7_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_7_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_7_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_7_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_7_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_7_io_pSumOut_bits),
    .io_stateOut(pes_2_7_io_stateOut)
  );
  dataSwitch dss_2_7 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_7_io_dataIn_ready),
    .io_dataIn_valid(dss_2_7_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_7_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_7_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_7_io_filter_ready),
    .io_filter_valid(dss_2_7_io_filter_valid),
    .io_filter_bits(dss_2_7_io_filter_bits),
    .io_ifmap_ready(dss_2_7_io_ifmap_ready),
    .io_ifmap_valid(dss_2_7_io_ifmap_valid),
    .io_ifmap_bits(dss_2_7_io_ifmap_bits),
    .io_pSum_ready(dss_2_7_io_pSum_ready),
    .io_pSum_valid(dss_2_7_io_pSum_valid),
    .io_pSum_bits(dss_2_7_io_pSum_bits)
  );
  Node_59 NoC_2_9 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_9_clock),
    .reset(NoC_2_9_reset),
    .io_dataPackageIn_ready(NoC_2_9_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_9_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_9_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_9_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_9_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_9_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_9_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_9_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_9_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_8 ( // @[PEArray.scala 36:24]
    .clock(pes_2_8_clock),
    .reset(pes_2_8_reset),
    .io_stateSW(pes_2_8_io_stateSW),
    .io_peconfig_ready(pes_2_8_io_peconfig_ready),
    .io_peconfig_valid(pes_2_8_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_8_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_8_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_8_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_8_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_8_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_8_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_8_io_filter_ready),
    .io_filter_valid(pes_2_8_io_filter_valid),
    .io_filter_bits(pes_2_8_io_filter_bits),
    .io_ifmap_ready(pes_2_8_io_ifmap_ready),
    .io_ifmap_valid(pes_2_8_io_ifmap_valid),
    .io_ifmap_bits(pes_2_8_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_8_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_8_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_8_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_8_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_8_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_8_io_pSumOut_bits),
    .io_stateOut(pes_2_8_io_stateOut)
  );
  dataSwitch dss_2_8 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_8_io_dataIn_ready),
    .io_dataIn_valid(dss_2_8_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_8_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_8_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_8_io_filter_ready),
    .io_filter_valid(dss_2_8_io_filter_valid),
    .io_filter_bits(dss_2_8_io_filter_bits),
    .io_ifmap_ready(dss_2_8_io_ifmap_ready),
    .io_ifmap_valid(dss_2_8_io_ifmap_valid),
    .io_ifmap_bits(dss_2_8_io_ifmap_bits),
    .io_pSum_ready(dss_2_8_io_pSum_ready),
    .io_pSum_valid(dss_2_8_io_pSum_valid),
    .io_pSum_bits(dss_2_8_io_pSum_bits)
  );
  Node_60 NoC_2_10 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_10_clock),
    .reset(NoC_2_10_reset),
    .io_dataPackageIn_ready(NoC_2_10_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_10_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_10_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_10_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_10_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_10_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_10_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_10_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_10_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_9 ( // @[PEArray.scala 36:24]
    .clock(pes_2_9_clock),
    .reset(pes_2_9_reset),
    .io_stateSW(pes_2_9_io_stateSW),
    .io_peconfig_ready(pes_2_9_io_peconfig_ready),
    .io_peconfig_valid(pes_2_9_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_9_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_9_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_9_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_9_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_9_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_9_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_9_io_filter_ready),
    .io_filter_valid(pes_2_9_io_filter_valid),
    .io_filter_bits(pes_2_9_io_filter_bits),
    .io_ifmap_ready(pes_2_9_io_ifmap_ready),
    .io_ifmap_valid(pes_2_9_io_ifmap_valid),
    .io_ifmap_bits(pes_2_9_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_9_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_9_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_9_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_9_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_9_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_9_io_pSumOut_bits),
    .io_stateOut(pes_2_9_io_stateOut)
  );
  dataSwitch dss_2_9 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_9_io_dataIn_ready),
    .io_dataIn_valid(dss_2_9_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_9_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_9_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_9_io_filter_ready),
    .io_filter_valid(dss_2_9_io_filter_valid),
    .io_filter_bits(dss_2_9_io_filter_bits),
    .io_ifmap_ready(dss_2_9_io_ifmap_ready),
    .io_ifmap_valid(dss_2_9_io_ifmap_valid),
    .io_ifmap_bits(dss_2_9_io_ifmap_bits),
    .io_pSum_ready(dss_2_9_io_pSum_ready),
    .io_pSum_valid(dss_2_9_io_pSum_valid),
    .io_pSum_bits(dss_2_9_io_pSum_bits)
  );
  Node_61 NoC_2_11 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_11_clock),
    .reset(NoC_2_11_reset),
    .io_dataPackageIn_ready(NoC_2_11_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_11_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_11_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_11_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_11_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_11_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_11_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_11_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_11_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_10 ( // @[PEArray.scala 36:24]
    .clock(pes_2_10_clock),
    .reset(pes_2_10_reset),
    .io_stateSW(pes_2_10_io_stateSW),
    .io_peconfig_ready(pes_2_10_io_peconfig_ready),
    .io_peconfig_valid(pes_2_10_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_10_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_10_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_10_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_10_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_10_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_10_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_10_io_filter_ready),
    .io_filter_valid(pes_2_10_io_filter_valid),
    .io_filter_bits(pes_2_10_io_filter_bits),
    .io_ifmap_ready(pes_2_10_io_ifmap_ready),
    .io_ifmap_valid(pes_2_10_io_ifmap_valid),
    .io_ifmap_bits(pes_2_10_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_10_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_10_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_10_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_10_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_10_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_10_io_pSumOut_bits),
    .io_stateOut(pes_2_10_io_stateOut)
  );
  dataSwitch dss_2_10 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_10_io_dataIn_ready),
    .io_dataIn_valid(dss_2_10_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_10_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_10_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_10_io_filter_ready),
    .io_filter_valid(dss_2_10_io_filter_valid),
    .io_filter_bits(dss_2_10_io_filter_bits),
    .io_ifmap_ready(dss_2_10_io_ifmap_ready),
    .io_ifmap_valid(dss_2_10_io_ifmap_valid),
    .io_ifmap_bits(dss_2_10_io_ifmap_bits),
    .io_pSum_ready(dss_2_10_io_pSum_ready),
    .io_pSum_valid(dss_2_10_io_pSum_valid),
    .io_pSum_bits(dss_2_10_io_pSum_bits)
  );
  Node_62 NoC_2_12 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_12_clock),
    .reset(NoC_2_12_reset),
    .io_dataPackageIn_ready(NoC_2_12_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_12_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_12_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_12_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_12_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_12_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_12_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_12_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_12_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_11 ( // @[PEArray.scala 36:24]
    .clock(pes_2_11_clock),
    .reset(pes_2_11_reset),
    .io_stateSW(pes_2_11_io_stateSW),
    .io_peconfig_ready(pes_2_11_io_peconfig_ready),
    .io_peconfig_valid(pes_2_11_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_11_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_11_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_11_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_11_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_11_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_11_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_11_io_filter_ready),
    .io_filter_valid(pes_2_11_io_filter_valid),
    .io_filter_bits(pes_2_11_io_filter_bits),
    .io_ifmap_ready(pes_2_11_io_ifmap_ready),
    .io_ifmap_valid(pes_2_11_io_ifmap_valid),
    .io_ifmap_bits(pes_2_11_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_11_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_11_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_11_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_11_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_11_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_11_io_pSumOut_bits),
    .io_stateOut(pes_2_11_io_stateOut)
  );
  dataSwitch dss_2_11 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_11_io_dataIn_ready),
    .io_dataIn_valid(dss_2_11_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_11_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_11_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_11_io_filter_ready),
    .io_filter_valid(dss_2_11_io_filter_valid),
    .io_filter_bits(dss_2_11_io_filter_bits),
    .io_ifmap_ready(dss_2_11_io_ifmap_ready),
    .io_ifmap_valid(dss_2_11_io_ifmap_valid),
    .io_ifmap_bits(dss_2_11_io_ifmap_bits),
    .io_pSum_ready(dss_2_11_io_pSum_ready),
    .io_pSum_valid(dss_2_11_io_pSum_valid),
    .io_pSum_bits(dss_2_11_io_pSum_bits)
  );
  Node_63 NoC_2_13 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_13_clock),
    .reset(NoC_2_13_reset),
    .io_dataPackageIn_ready(NoC_2_13_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_13_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_13_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_13_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_13_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_13_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_13_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_13_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_13_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_12 ( // @[PEArray.scala 36:24]
    .clock(pes_2_12_clock),
    .reset(pes_2_12_reset),
    .io_stateSW(pes_2_12_io_stateSW),
    .io_peconfig_ready(pes_2_12_io_peconfig_ready),
    .io_peconfig_valid(pes_2_12_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_12_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_12_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_12_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_12_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_12_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_12_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_12_io_filter_ready),
    .io_filter_valid(pes_2_12_io_filter_valid),
    .io_filter_bits(pes_2_12_io_filter_bits),
    .io_ifmap_ready(pes_2_12_io_ifmap_ready),
    .io_ifmap_valid(pes_2_12_io_ifmap_valid),
    .io_ifmap_bits(pes_2_12_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_12_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_12_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_12_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_12_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_12_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_12_io_pSumOut_bits),
    .io_stateOut(pes_2_12_io_stateOut)
  );
  dataSwitch dss_2_12 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_12_io_dataIn_ready),
    .io_dataIn_valid(dss_2_12_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_12_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_12_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_12_io_filter_ready),
    .io_filter_valid(dss_2_12_io_filter_valid),
    .io_filter_bits(dss_2_12_io_filter_bits),
    .io_ifmap_ready(dss_2_12_io_ifmap_ready),
    .io_ifmap_valid(dss_2_12_io_ifmap_valid),
    .io_ifmap_bits(dss_2_12_io_ifmap_bits),
    .io_pSum_ready(dss_2_12_io_pSum_ready),
    .io_pSum_valid(dss_2_12_io_pSum_valid),
    .io_pSum_bits(dss_2_12_io_pSum_bits)
  );
  Node_64 NoC_2_14 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_14_clock),
    .reset(NoC_2_14_reset),
    .io_dataPackageIn_ready(NoC_2_14_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_14_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_14_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_14_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_14_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_14_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_14_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_14_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_14_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_13 ( // @[PEArray.scala 36:24]
    .clock(pes_2_13_clock),
    .reset(pes_2_13_reset),
    .io_stateSW(pes_2_13_io_stateSW),
    .io_peconfig_ready(pes_2_13_io_peconfig_ready),
    .io_peconfig_valid(pes_2_13_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_13_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_13_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_13_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_13_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_13_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_13_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_13_io_filter_ready),
    .io_filter_valid(pes_2_13_io_filter_valid),
    .io_filter_bits(pes_2_13_io_filter_bits),
    .io_ifmap_ready(pes_2_13_io_ifmap_ready),
    .io_ifmap_valid(pes_2_13_io_ifmap_valid),
    .io_ifmap_bits(pes_2_13_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_13_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_13_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_13_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_13_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_13_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_13_io_pSumOut_bits),
    .io_stateOut(pes_2_13_io_stateOut)
  );
  dataSwitch dss_2_13 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_13_io_dataIn_ready),
    .io_dataIn_valid(dss_2_13_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_13_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_13_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_13_io_filter_ready),
    .io_filter_valid(dss_2_13_io_filter_valid),
    .io_filter_bits(dss_2_13_io_filter_bits),
    .io_ifmap_ready(dss_2_13_io_ifmap_ready),
    .io_ifmap_valid(dss_2_13_io_ifmap_valid),
    .io_ifmap_bits(dss_2_13_io_ifmap_bits),
    .io_pSum_ready(dss_2_13_io_pSum_ready),
    .io_pSum_valid(dss_2_13_io_pSum_valid),
    .io_pSum_bits(dss_2_13_io_pSum_bits)
  );
  Node_65 NoC_2_15 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_15_clock),
    .reset(NoC_2_15_reset),
    .io_dataPackageIn_ready(NoC_2_15_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_15_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_15_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_15_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_15_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_15_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_15_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_15_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_15_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_14 ( // @[PEArray.scala 36:24]
    .clock(pes_2_14_clock),
    .reset(pes_2_14_reset),
    .io_stateSW(pes_2_14_io_stateSW),
    .io_peconfig_ready(pes_2_14_io_peconfig_ready),
    .io_peconfig_valid(pes_2_14_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_14_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_14_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_14_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_14_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_14_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_14_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_14_io_filter_ready),
    .io_filter_valid(pes_2_14_io_filter_valid),
    .io_filter_bits(pes_2_14_io_filter_bits),
    .io_ifmap_ready(pes_2_14_io_ifmap_ready),
    .io_ifmap_valid(pes_2_14_io_ifmap_valid),
    .io_ifmap_bits(pes_2_14_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_14_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_14_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_14_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_14_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_14_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_14_io_pSumOut_bits),
    .io_stateOut(pes_2_14_io_stateOut)
  );
  dataSwitch dss_2_14 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_14_io_dataIn_ready),
    .io_dataIn_valid(dss_2_14_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_14_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_14_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_14_io_filter_ready),
    .io_filter_valid(dss_2_14_io_filter_valid),
    .io_filter_bits(dss_2_14_io_filter_bits),
    .io_ifmap_ready(dss_2_14_io_ifmap_ready),
    .io_ifmap_valid(dss_2_14_io_ifmap_valid),
    .io_ifmap_bits(dss_2_14_io_ifmap_bits),
    .io_pSum_ready(dss_2_14_io_pSum_ready),
    .io_pSum_valid(dss_2_14_io_pSum_valid),
    .io_pSum_bits(dss_2_14_io_pSum_bits)
  );
  Node_66 NoC_2_16 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_16_clock),
    .reset(NoC_2_16_reset),
    .io_dataPackageIn_ready(NoC_2_16_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_16_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_16_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_16_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_16_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_16_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_16_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_16_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_16_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_15 ( // @[PEArray.scala 36:24]
    .clock(pes_2_15_clock),
    .reset(pes_2_15_reset),
    .io_stateSW(pes_2_15_io_stateSW),
    .io_peconfig_ready(pes_2_15_io_peconfig_ready),
    .io_peconfig_valid(pes_2_15_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_15_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_15_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_15_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_15_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_15_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_15_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_15_io_filter_ready),
    .io_filter_valid(pes_2_15_io_filter_valid),
    .io_filter_bits(pes_2_15_io_filter_bits),
    .io_ifmap_ready(pes_2_15_io_ifmap_ready),
    .io_ifmap_valid(pes_2_15_io_ifmap_valid),
    .io_ifmap_bits(pes_2_15_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_15_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_15_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_15_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_15_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_15_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_15_io_pSumOut_bits),
    .io_stateOut(pes_2_15_io_stateOut)
  );
  dataSwitch dss_2_15 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_15_io_dataIn_ready),
    .io_dataIn_valid(dss_2_15_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_15_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_15_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_15_io_filter_ready),
    .io_filter_valid(dss_2_15_io_filter_valid),
    .io_filter_bits(dss_2_15_io_filter_bits),
    .io_ifmap_ready(dss_2_15_io_ifmap_ready),
    .io_ifmap_valid(dss_2_15_io_ifmap_valid),
    .io_ifmap_bits(dss_2_15_io_ifmap_bits),
    .io_pSum_ready(dss_2_15_io_pSum_ready),
    .io_pSum_valid(dss_2_15_io_pSum_valid),
    .io_pSum_bits(dss_2_15_io_pSum_bits)
  );
  Node_67 NoC_2_17 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_17_clock),
    .reset(NoC_2_17_reset),
    .io_dataPackageIn_ready(NoC_2_17_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_17_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_17_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_17_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_17_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_17_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_17_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_17_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_17_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_16 ( // @[PEArray.scala 36:24]
    .clock(pes_2_16_clock),
    .reset(pes_2_16_reset),
    .io_stateSW(pes_2_16_io_stateSW),
    .io_peconfig_ready(pes_2_16_io_peconfig_ready),
    .io_peconfig_valid(pes_2_16_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_16_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_16_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_16_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_16_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_16_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_16_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_16_io_filter_ready),
    .io_filter_valid(pes_2_16_io_filter_valid),
    .io_filter_bits(pes_2_16_io_filter_bits),
    .io_ifmap_ready(pes_2_16_io_ifmap_ready),
    .io_ifmap_valid(pes_2_16_io_ifmap_valid),
    .io_ifmap_bits(pes_2_16_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_16_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_16_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_16_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_16_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_16_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_16_io_pSumOut_bits),
    .io_stateOut(pes_2_16_io_stateOut)
  );
  dataSwitch dss_2_16 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_16_io_dataIn_ready),
    .io_dataIn_valid(dss_2_16_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_16_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_16_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_16_io_filter_ready),
    .io_filter_valid(dss_2_16_io_filter_valid),
    .io_filter_bits(dss_2_16_io_filter_bits),
    .io_ifmap_ready(dss_2_16_io_ifmap_ready),
    .io_ifmap_valid(dss_2_16_io_ifmap_valid),
    .io_ifmap_bits(dss_2_16_io_ifmap_bits),
    .io_pSum_ready(dss_2_16_io_pSum_ready),
    .io_pSum_valid(dss_2_16_io_pSum_valid),
    .io_pSum_bits(dss_2_16_io_pSum_bits)
  );
  Node_68 NoC_2_18 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_18_clock),
    .reset(NoC_2_18_reset),
    .io_dataPackageIn_ready(NoC_2_18_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_18_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_18_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_18_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_18_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_18_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_18_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_18_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_18_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_17 ( // @[PEArray.scala 36:24]
    .clock(pes_2_17_clock),
    .reset(pes_2_17_reset),
    .io_stateSW(pes_2_17_io_stateSW),
    .io_peconfig_ready(pes_2_17_io_peconfig_ready),
    .io_peconfig_valid(pes_2_17_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_17_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_17_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_17_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_17_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_17_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_17_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_17_io_filter_ready),
    .io_filter_valid(pes_2_17_io_filter_valid),
    .io_filter_bits(pes_2_17_io_filter_bits),
    .io_ifmap_ready(pes_2_17_io_ifmap_ready),
    .io_ifmap_valid(pes_2_17_io_ifmap_valid),
    .io_ifmap_bits(pes_2_17_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_17_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_17_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_17_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_17_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_17_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_17_io_pSumOut_bits),
    .io_stateOut(pes_2_17_io_stateOut)
  );
  dataSwitch dss_2_17 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_17_io_dataIn_ready),
    .io_dataIn_valid(dss_2_17_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_17_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_17_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_17_io_filter_ready),
    .io_filter_valid(dss_2_17_io_filter_valid),
    .io_filter_bits(dss_2_17_io_filter_bits),
    .io_ifmap_ready(dss_2_17_io_ifmap_ready),
    .io_ifmap_valid(dss_2_17_io_ifmap_valid),
    .io_ifmap_bits(dss_2_17_io_ifmap_bits),
    .io_pSum_ready(dss_2_17_io_pSum_ready),
    .io_pSum_valid(dss_2_17_io_pSum_valid),
    .io_pSum_bits(dss_2_17_io_pSum_bits)
  );
  Node_69 NoC_2_19 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_19_clock),
    .reset(NoC_2_19_reset),
    .io_dataPackageIn_ready(NoC_2_19_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_19_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_19_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_19_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_19_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_19_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_19_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_19_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_19_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_18 ( // @[PEArray.scala 36:24]
    .clock(pes_2_18_clock),
    .reset(pes_2_18_reset),
    .io_stateSW(pes_2_18_io_stateSW),
    .io_peconfig_ready(pes_2_18_io_peconfig_ready),
    .io_peconfig_valid(pes_2_18_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_18_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_18_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_18_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_18_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_18_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_18_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_18_io_filter_ready),
    .io_filter_valid(pes_2_18_io_filter_valid),
    .io_filter_bits(pes_2_18_io_filter_bits),
    .io_ifmap_ready(pes_2_18_io_ifmap_ready),
    .io_ifmap_valid(pes_2_18_io_ifmap_valid),
    .io_ifmap_bits(pes_2_18_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_18_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_18_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_18_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_18_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_18_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_18_io_pSumOut_bits),
    .io_stateOut(pes_2_18_io_stateOut)
  );
  dataSwitch dss_2_18 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_18_io_dataIn_ready),
    .io_dataIn_valid(dss_2_18_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_18_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_18_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_18_io_filter_ready),
    .io_filter_valid(dss_2_18_io_filter_valid),
    .io_filter_bits(dss_2_18_io_filter_bits),
    .io_ifmap_ready(dss_2_18_io_ifmap_ready),
    .io_ifmap_valid(dss_2_18_io_ifmap_valid),
    .io_ifmap_bits(dss_2_18_io_ifmap_bits),
    .io_pSum_ready(dss_2_18_io_pSum_ready),
    .io_pSum_valid(dss_2_18_io_pSum_valid),
    .io_pSum_bits(dss_2_18_io_pSum_bits)
  );
  Node_70 NoC_2_20 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_20_clock),
    .reset(NoC_2_20_reset),
    .io_dataPackageIn_ready(NoC_2_20_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_20_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_20_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_20_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_20_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_20_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_20_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_20_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_20_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_19 ( // @[PEArray.scala 36:24]
    .clock(pes_2_19_clock),
    .reset(pes_2_19_reset),
    .io_stateSW(pes_2_19_io_stateSW),
    .io_peconfig_ready(pes_2_19_io_peconfig_ready),
    .io_peconfig_valid(pes_2_19_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_19_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_19_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_19_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_19_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_19_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_19_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_19_io_filter_ready),
    .io_filter_valid(pes_2_19_io_filter_valid),
    .io_filter_bits(pes_2_19_io_filter_bits),
    .io_ifmap_ready(pes_2_19_io_ifmap_ready),
    .io_ifmap_valid(pes_2_19_io_ifmap_valid),
    .io_ifmap_bits(pes_2_19_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_19_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_19_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_19_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_19_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_19_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_19_io_pSumOut_bits),
    .io_stateOut(pes_2_19_io_stateOut)
  );
  dataSwitch dss_2_19 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_19_io_dataIn_ready),
    .io_dataIn_valid(dss_2_19_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_19_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_19_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_19_io_filter_ready),
    .io_filter_valid(dss_2_19_io_filter_valid),
    .io_filter_bits(dss_2_19_io_filter_bits),
    .io_ifmap_ready(dss_2_19_io_ifmap_ready),
    .io_ifmap_valid(dss_2_19_io_ifmap_valid),
    .io_ifmap_bits(dss_2_19_io_ifmap_bits),
    .io_pSum_ready(dss_2_19_io_pSum_ready),
    .io_pSum_valid(dss_2_19_io_pSum_valid),
    .io_pSum_bits(dss_2_19_io_pSum_bits)
  );
  Node_71 NoC_2_21 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_21_clock),
    .reset(NoC_2_21_reset),
    .io_dataPackageIn_ready(NoC_2_21_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_21_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_21_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_21_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_21_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_21_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_21_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_21_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_21_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_20 ( // @[PEArray.scala 36:24]
    .clock(pes_2_20_clock),
    .reset(pes_2_20_reset),
    .io_stateSW(pes_2_20_io_stateSW),
    .io_peconfig_ready(pes_2_20_io_peconfig_ready),
    .io_peconfig_valid(pes_2_20_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_20_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_20_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_20_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_20_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_20_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_20_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_20_io_filter_ready),
    .io_filter_valid(pes_2_20_io_filter_valid),
    .io_filter_bits(pes_2_20_io_filter_bits),
    .io_ifmap_ready(pes_2_20_io_ifmap_ready),
    .io_ifmap_valid(pes_2_20_io_ifmap_valid),
    .io_ifmap_bits(pes_2_20_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_20_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_20_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_20_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_20_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_20_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_20_io_pSumOut_bits),
    .io_stateOut(pes_2_20_io_stateOut)
  );
  dataSwitch dss_2_20 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_20_io_dataIn_ready),
    .io_dataIn_valid(dss_2_20_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_20_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_20_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_20_io_filter_ready),
    .io_filter_valid(dss_2_20_io_filter_valid),
    .io_filter_bits(dss_2_20_io_filter_bits),
    .io_ifmap_ready(dss_2_20_io_ifmap_ready),
    .io_ifmap_valid(dss_2_20_io_ifmap_valid),
    .io_ifmap_bits(dss_2_20_io_ifmap_bits),
    .io_pSum_ready(dss_2_20_io_pSum_ready),
    .io_pSum_valid(dss_2_20_io_pSum_valid),
    .io_pSum_bits(dss_2_20_io_pSum_bits)
  );
  Node_72 NoC_2_22 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_22_clock),
    .reset(NoC_2_22_reset),
    .io_dataPackageIn_ready(NoC_2_22_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_22_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_22_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_22_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_22_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_22_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_22_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_22_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_22_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_21 ( // @[PEArray.scala 36:24]
    .clock(pes_2_21_clock),
    .reset(pes_2_21_reset),
    .io_stateSW(pes_2_21_io_stateSW),
    .io_peconfig_ready(pes_2_21_io_peconfig_ready),
    .io_peconfig_valid(pes_2_21_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_21_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_21_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_21_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_21_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_21_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_21_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_21_io_filter_ready),
    .io_filter_valid(pes_2_21_io_filter_valid),
    .io_filter_bits(pes_2_21_io_filter_bits),
    .io_ifmap_ready(pes_2_21_io_ifmap_ready),
    .io_ifmap_valid(pes_2_21_io_ifmap_valid),
    .io_ifmap_bits(pes_2_21_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_21_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_21_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_21_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_21_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_21_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_21_io_pSumOut_bits),
    .io_stateOut(pes_2_21_io_stateOut)
  );
  dataSwitch dss_2_21 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_21_io_dataIn_ready),
    .io_dataIn_valid(dss_2_21_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_21_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_21_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_21_io_filter_ready),
    .io_filter_valid(dss_2_21_io_filter_valid),
    .io_filter_bits(dss_2_21_io_filter_bits),
    .io_ifmap_ready(dss_2_21_io_ifmap_ready),
    .io_ifmap_valid(dss_2_21_io_ifmap_valid),
    .io_ifmap_bits(dss_2_21_io_ifmap_bits),
    .io_pSum_ready(dss_2_21_io_pSum_ready),
    .io_pSum_valid(dss_2_21_io_pSum_valid),
    .io_pSum_bits(dss_2_21_io_pSum_bits)
  );
  Node_73 NoC_2_23 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_23_clock),
    .reset(NoC_2_23_reset),
    .io_dataPackageIn_ready(NoC_2_23_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_23_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_23_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_23_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_23_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_23_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_23_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_23_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_23_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_22 ( // @[PEArray.scala 36:24]
    .clock(pes_2_22_clock),
    .reset(pes_2_22_reset),
    .io_stateSW(pes_2_22_io_stateSW),
    .io_peconfig_ready(pes_2_22_io_peconfig_ready),
    .io_peconfig_valid(pes_2_22_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_22_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_22_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_22_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_22_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_22_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_22_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_22_io_filter_ready),
    .io_filter_valid(pes_2_22_io_filter_valid),
    .io_filter_bits(pes_2_22_io_filter_bits),
    .io_ifmap_ready(pes_2_22_io_ifmap_ready),
    .io_ifmap_valid(pes_2_22_io_ifmap_valid),
    .io_ifmap_bits(pes_2_22_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_22_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_22_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_22_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_22_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_22_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_22_io_pSumOut_bits),
    .io_stateOut(pes_2_22_io_stateOut)
  );
  dataSwitch dss_2_22 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_22_io_dataIn_ready),
    .io_dataIn_valid(dss_2_22_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_22_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_22_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_22_io_filter_ready),
    .io_filter_valid(dss_2_22_io_filter_valid),
    .io_filter_bits(dss_2_22_io_filter_bits),
    .io_ifmap_ready(dss_2_22_io_ifmap_ready),
    .io_ifmap_valid(dss_2_22_io_ifmap_valid),
    .io_ifmap_bits(dss_2_22_io_ifmap_bits),
    .io_pSum_ready(dss_2_22_io_pSum_ready),
    .io_pSum_valid(dss_2_22_io_pSum_valid),
    .io_pSum_bits(dss_2_22_io_pSum_bits)
  );
  Node_74 NoC_2_24 ( // @[PEArray.scala 34:24]
    .clock(NoC_2_24_clock),
    .reset(NoC_2_24_reset),
    .io_dataPackageIn_ready(NoC_2_24_io_dataPackageIn_ready),
    .io_dataPackageIn_valid(NoC_2_24_io_dataPackageIn_valid),
    .io_dataPackageIn_bits_data(NoC_2_24_io_dataPackageIn_bits_data),
    .io_dataPackageIn_bits_dataType(NoC_2_24_io_dataPackageIn_bits_dataType),
    .io_dataPackageIn_bits_positon_col(NoC_2_24_io_dataPackageIn_bits_positon_col),
    .io_dataPackageOut_ready(NoC_2_24_io_dataPackageOut_ready),
    .io_dataPackageOut_valid(NoC_2_24_io_dataPackageOut_valid),
    .io_dataPackageOut_bits_data(NoC_2_24_io_dataPackageOut_bits_data),
    .io_dataPackageOut_bits_dataType(NoC_2_24_io_dataPackageOut_bits_dataType)
  );
  PETop pes_2_23 ( // @[PEArray.scala 36:24]
    .clock(pes_2_23_clock),
    .reset(pes_2_23_reset),
    .io_stateSW(pes_2_23_io_stateSW),
    .io_peconfig_ready(pes_2_23_io_peconfig_ready),
    .io_peconfig_valid(pes_2_23_io_peconfig_valid),
    .io_peconfig_bits_ichannelNum(pes_2_23_io_peconfig_bits_ichannelNum),
    .io_peconfig_bits_ochannelNum(pes_2_23_io_peconfig_bits_ochannelNum),
    .io_peconfig_bits_ofmapW(pes_2_23_io_peconfig_bits_ofmapW),
    .io_peconfig_bits_stepW(pes_2_23_io_peconfig_bits_stepW),
    .io_peconfig_bits_filterLen(pes_2_23_io_peconfig_bits_filterLen),
    .io_peconfig_bits_ifmapLen(pes_2_23_io_peconfig_bits_ifmapLen),
    .io_filter_ready(pes_2_23_io_filter_ready),
    .io_filter_valid(pes_2_23_io_filter_valid),
    .io_filter_bits(pes_2_23_io_filter_bits),
    .io_ifmap_ready(pes_2_23_io_ifmap_ready),
    .io_ifmap_valid(pes_2_23_io_ifmap_valid),
    .io_ifmap_bits(pes_2_23_io_ifmap_bits),
    .io_pSumIn_ready(pes_2_23_io_pSumIn_ready),
    .io_pSumIn_valid(pes_2_23_io_pSumIn_valid),
    .io_pSumIn_bits(pes_2_23_io_pSumIn_bits),
    .io_pSumOut_ready(pes_2_23_io_pSumOut_ready),
    .io_pSumOut_valid(pes_2_23_io_pSumOut_valid),
    .io_pSumOut_bits(pes_2_23_io_pSumOut_bits),
    .io_stateOut(pes_2_23_io_stateOut)
  );
  dataSwitch dss_2_23 ( // @[PEArray.scala 37:24]
    .io_dataIn_ready(dss_2_23_io_dataIn_ready),
    .io_dataIn_valid(dss_2_23_io_dataIn_valid),
    .io_dataIn_bits_data(dss_2_23_io_dataIn_bits_data),
    .io_dataIn_bits_dataType(dss_2_23_io_dataIn_bits_dataType),
    .io_filter_ready(dss_2_23_io_filter_ready),
    .io_filter_valid(dss_2_23_io_filter_valid),
    .io_filter_bits(dss_2_23_io_filter_bits),
    .io_ifmap_ready(dss_2_23_io_ifmap_ready),
    .io_ifmap_valid(dss_2_23_io_ifmap_valid),
    .io_ifmap_bits(dss_2_23_io_ifmap_bits),
    .io_pSum_ready(dss_2_23_io_pSum_ready),
    .io_pSum_valid(dss_2_23_io_pSum_valid),
    .io_pSum_bits(dss_2_23_io_pSum_bits)
  );
  assign io_dataIn_ready = NoC_0_0_io_dataPackageIn_ready | NoC_1_0_io_dataPackageIn_ready |
    NoC_2_0_io_dataPackageIn_ready; // @[PEArray.scala 87:70]
  assign io_peconfig_ready = _T_250 | pes_2_13_io_peconfig_ready | pes_2_14_io_peconfig_ready |
    pes_2_15_io_peconfig_ready | pes_2_16_io_peconfig_ready | pes_2_17_io_peconfig_ready | pes_2_18_io_peconfig_ready |
    pes_2_19_io_peconfig_ready | pes_2_20_io_peconfig_ready | pes_2_21_io_peconfig_ready | pes_2_22_io_peconfig_ready |
    pes_2_23_io_peconfig_ready; // @[PEArray.scala 106:77]
  assign io_oSumOut_0_valid = pes_2_0_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_0_bits = configReg_relu & $signed(pes_2_0_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_0_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_1_valid = pes_2_1_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_1_bits = configReg_relu & $signed(pes_2_1_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_1_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_2_valid = pes_2_2_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_2_bits = configReg_relu & $signed(pes_2_2_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_2_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_3_valid = pes_2_3_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_3_bits = configReg_relu & $signed(pes_2_3_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_3_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_4_valid = pes_2_4_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_4_bits = configReg_relu & $signed(pes_2_4_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_4_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_5_valid = pes_2_5_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_5_bits = configReg_relu & $signed(pes_2_5_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_5_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_6_valid = pes_2_6_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_6_bits = configReg_relu & $signed(pes_2_6_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_6_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_7_valid = pes_2_7_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_7_bits = configReg_relu & $signed(pes_2_7_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_7_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_8_valid = pes_2_8_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_8_bits = configReg_relu & $signed(pes_2_8_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_8_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_9_valid = pes_2_9_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_9_bits = configReg_relu & $signed(pes_2_9_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_9_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_10_valid = pes_2_10_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_10_bits = configReg_relu & $signed(pes_2_10_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_10_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_11_valid = pes_2_11_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_11_bits = configReg_relu & $signed(pes_2_11_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_11_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_12_valid = pes_2_12_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_12_bits = configReg_relu & $signed(pes_2_12_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_12_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_13_valid = pes_2_13_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_13_bits = configReg_relu & $signed(pes_2_13_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_13_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_14_valid = pes_2_14_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_14_bits = configReg_relu & $signed(pes_2_14_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_14_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_15_valid = pes_2_15_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_15_bits = configReg_relu & $signed(pes_2_15_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_15_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_16_valid = pes_2_16_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_16_bits = configReg_relu & $signed(pes_2_16_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_16_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_17_valid = pes_2_17_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_17_bits = configReg_relu & $signed(pes_2_17_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_17_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_18_valid = pes_2_18_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_18_bits = configReg_relu & $signed(pes_2_18_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_18_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_19_valid = pes_2_19_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_19_bits = configReg_relu & $signed(pes_2_19_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_19_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_20_valid = pes_2_20_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_20_bits = configReg_relu & $signed(pes_2_20_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_20_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_21_valid = pes_2_21_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_21_bits = configReg_relu & $signed(pes_2_21_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_21_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_22_valid = pes_2_22_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_22_bits = configReg_relu & $signed(pes_2_22_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_22_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_oSumOut_23_valid = pes_2_23_io_pSumOut_valid; // @[PEArray.scala 52:33]
  assign io_oSumOut_23_bits = configReg_relu & $signed(pes_2_23_io_pSumOut_bits) < 20'sh0 ? $signed(20'sh0) : $signed(
    pes_2_23_io_pSumOut_bits); // @[PEArray.scala 55:67 PEArray.scala 56:34 PEArray.scala 58:34]
  assign io_done = doneReg; // @[PEArray.scala 18:11]
  assign NoC_0_0_clock = clock;
  assign NoC_0_0_reset = reset;
  assign NoC_0_0_io_dataPackageIn_valid = io_dataIn_valid; // @[PEArray.scala 84:35]
  assign NoC_0_0_io_dataPackageIn_bits_data = io_dataIn_bits_data; // @[PEArray.scala 85:34]
  assign NoC_0_0_io_dataPackageIn_bits_dataType = io_dataIn_bits_dataType; // @[PEArray.scala 85:34]
  assign NoC_0_0_io_dataPackageIn_bits_positon_row = io_dataIn_bits_positon_row; // @[PEArray.scala 85:34]
  assign NoC_0_0_io_dataPackageIn_bits_positon_col = io_dataIn_bits_positon_col; // @[PEArray.scala 85:34]
  assign NoC_0_0_io_dataPackageOut_ready = NoC_0_1_io_dataPackageIn_ready | NoC_0_2_io_dataPackageIn_ready |
    NoC_0_3_io_dataPackageIn_ready | NoC_0_4_io_dataPackageIn_ready | NoC_0_5_io_dataPackageIn_ready |
    NoC_0_6_io_dataPackageIn_ready | NoC_0_7_io_dataPackageIn_ready | NoC_0_8_io_dataPackageIn_ready |
    NoC_0_9_io_dataPackageIn_ready | NoC_0_10_io_dataPackageIn_ready | NoC_0_11_io_dataPackageIn_ready |
    NoC_0_12_io_dataPackageIn_ready | NoC_0_13_io_dataPackageIn_ready | NoC_0_14_io_dataPackageIn_ready |
    NoC_0_15_io_dataPackageIn_ready | NoC_0_16_io_dataPackageIn_ready | NoC_0_17_io_dataPackageIn_ready |
    NoC_0_18_io_dataPackageIn_ready | NoC_0_19_io_dataPackageIn_ready | NoC_0_20_io_dataPackageIn_ready |
    NoC_0_21_io_dataPackageIn_ready | NoC_0_22_io_dataPackageIn_ready | NoC_0_23_io_dataPackageIn_ready |
    NoC_0_24_io_dataPackageIn_ready; // @[PEArray.scala 83:17]
  assign NoC_0_1_clock = clock;
  assign NoC_0_1_reset = reset;
  assign NoC_0_1_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_1_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_1_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_1_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_1_io_dataPackageOut_ready = dss_0_0_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_0_clock = clock;
  assign pes_0_0_reset = reset;
  assign pes_0_0_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_0_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_0_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_0_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_0_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_0_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_0_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_0_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_0_io_filter_valid = dss_0_0_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_0_io_filter_bits = dss_0_0_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_0_io_ifmap_valid = dss_0_0_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_0_io_ifmap_bits = dss_0_0_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_0_io_pSumIn_valid = dss_0_0_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_0_io_pSumIn_bits = {{4{dss_0_0_io_pSum_bits[15]}},dss_0_0_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_0_io_pSumOut_ready = pes_1_0_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_0_io_dataIn_valid = NoC_0_1_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_0_io_dataIn_bits_data = {{11{NoC_0_1_io_dataPackageOut_bits_data[4]}},NoC_0_1_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_0_0_io_dataIn_bits_dataType = NoC_0_1_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_0_io_filter_ready = pes_0_0_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_0_io_ifmap_ready = pes_0_0_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_0_io_pSum_ready = pes_0_0_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_2_clock = clock;
  assign NoC_0_2_reset = reset;
  assign NoC_0_2_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_2_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_2_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_2_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_2_io_dataPackageOut_ready = dss_0_1_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_1_clock = clock;
  assign pes_0_1_reset = reset;
  assign pes_0_1_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_1_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_1_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_1_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_1_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_1_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_1_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_1_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_1_io_filter_valid = dss_0_1_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_1_io_filter_bits = dss_0_1_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_1_io_ifmap_valid = dss_0_1_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_1_io_ifmap_bits = dss_0_1_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_1_io_pSumIn_valid = dss_0_1_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_1_io_pSumIn_bits = {{4{dss_0_1_io_pSum_bits[15]}},dss_0_1_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_1_io_pSumOut_ready = pes_1_1_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_1_io_dataIn_valid = NoC_0_2_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_1_io_dataIn_bits_data = {{11{NoC_0_2_io_dataPackageOut_bits_data[4]}},NoC_0_2_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_0_1_io_dataIn_bits_dataType = NoC_0_2_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_1_io_filter_ready = pes_0_1_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_1_io_ifmap_ready = pes_0_1_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_1_io_pSum_ready = pes_0_1_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_3_clock = clock;
  assign NoC_0_3_reset = reset;
  assign NoC_0_3_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_3_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_3_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_3_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_3_io_dataPackageOut_ready = dss_0_2_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_2_clock = clock;
  assign pes_0_2_reset = reset;
  assign pes_0_2_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_2_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_2_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_2_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_2_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_2_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_2_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_2_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_2_io_filter_valid = dss_0_2_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_2_io_filter_bits = dss_0_2_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_2_io_ifmap_valid = dss_0_2_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_2_io_ifmap_bits = dss_0_2_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_2_io_pSumIn_valid = dss_0_2_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_2_io_pSumIn_bits = {{4{dss_0_2_io_pSum_bits[15]}},dss_0_2_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_2_io_pSumOut_ready = pes_1_2_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_2_io_dataIn_valid = NoC_0_3_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_2_io_dataIn_bits_data = {{11{NoC_0_3_io_dataPackageOut_bits_data[4]}},NoC_0_3_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_0_2_io_dataIn_bits_dataType = NoC_0_3_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_2_io_filter_ready = pes_0_2_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_2_io_ifmap_ready = pes_0_2_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_2_io_pSum_ready = pes_0_2_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_4_clock = clock;
  assign NoC_0_4_reset = reset;
  assign NoC_0_4_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_4_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_4_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_4_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_4_io_dataPackageOut_ready = dss_0_3_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_3_clock = clock;
  assign pes_0_3_reset = reset;
  assign pes_0_3_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_3_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_3_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_3_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_3_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_3_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_3_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_3_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_3_io_filter_valid = dss_0_3_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_3_io_filter_bits = dss_0_3_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_3_io_ifmap_valid = dss_0_3_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_3_io_ifmap_bits = dss_0_3_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_3_io_pSumIn_valid = dss_0_3_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_3_io_pSumIn_bits = {{4{dss_0_3_io_pSum_bits[15]}},dss_0_3_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_3_io_pSumOut_ready = pes_1_3_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_3_io_dataIn_valid = NoC_0_4_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_3_io_dataIn_bits_data = {{11{NoC_0_4_io_dataPackageOut_bits_data[4]}},NoC_0_4_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_0_3_io_dataIn_bits_dataType = NoC_0_4_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_3_io_filter_ready = pes_0_3_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_3_io_ifmap_ready = pes_0_3_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_3_io_pSum_ready = pes_0_3_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_5_clock = clock;
  assign NoC_0_5_reset = reset;
  assign NoC_0_5_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_5_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_5_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_5_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_5_io_dataPackageOut_ready = dss_0_4_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_4_clock = clock;
  assign pes_0_4_reset = reset;
  assign pes_0_4_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_4_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_4_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_4_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_4_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_4_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_4_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_4_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_4_io_filter_valid = dss_0_4_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_4_io_filter_bits = dss_0_4_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_4_io_ifmap_valid = dss_0_4_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_4_io_ifmap_bits = dss_0_4_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_4_io_pSumIn_valid = dss_0_4_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_4_io_pSumIn_bits = {{4{dss_0_4_io_pSum_bits[15]}},dss_0_4_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_4_io_pSumOut_ready = pes_1_4_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_4_io_dataIn_valid = NoC_0_5_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_4_io_dataIn_bits_data = {{11{NoC_0_5_io_dataPackageOut_bits_data[4]}},NoC_0_5_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_0_4_io_dataIn_bits_dataType = NoC_0_5_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_4_io_filter_ready = pes_0_4_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_4_io_ifmap_ready = pes_0_4_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_4_io_pSum_ready = pes_0_4_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_6_clock = clock;
  assign NoC_0_6_reset = reset;
  assign NoC_0_6_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_6_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_6_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_6_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_6_io_dataPackageOut_ready = dss_0_5_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_5_clock = clock;
  assign pes_0_5_reset = reset;
  assign pes_0_5_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_5_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_5_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_5_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_5_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_5_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_5_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_5_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_5_io_filter_valid = dss_0_5_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_5_io_filter_bits = dss_0_5_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_5_io_ifmap_valid = dss_0_5_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_5_io_ifmap_bits = dss_0_5_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_5_io_pSumIn_valid = dss_0_5_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_5_io_pSumIn_bits = {{4{dss_0_5_io_pSum_bits[15]}},dss_0_5_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_5_io_pSumOut_ready = pes_1_5_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_5_io_dataIn_valid = NoC_0_6_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_5_io_dataIn_bits_data = {{11{NoC_0_6_io_dataPackageOut_bits_data[4]}},NoC_0_6_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_0_5_io_dataIn_bits_dataType = NoC_0_6_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_5_io_filter_ready = pes_0_5_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_5_io_ifmap_ready = pes_0_5_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_5_io_pSum_ready = pes_0_5_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_7_clock = clock;
  assign NoC_0_7_reset = reset;
  assign NoC_0_7_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_7_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_7_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_7_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_7_io_dataPackageOut_ready = dss_0_6_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_6_clock = clock;
  assign pes_0_6_reset = reset;
  assign pes_0_6_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_6_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_6_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_6_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_6_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_6_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_6_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_6_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_6_io_filter_valid = dss_0_6_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_6_io_filter_bits = dss_0_6_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_6_io_ifmap_valid = dss_0_6_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_6_io_ifmap_bits = dss_0_6_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_6_io_pSumIn_valid = dss_0_6_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_6_io_pSumIn_bits = {{4{dss_0_6_io_pSum_bits[15]}},dss_0_6_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_6_io_pSumOut_ready = pes_1_6_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_6_io_dataIn_valid = NoC_0_7_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_6_io_dataIn_bits_data = {{11{NoC_0_7_io_dataPackageOut_bits_data[4]}},NoC_0_7_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_0_6_io_dataIn_bits_dataType = NoC_0_7_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_6_io_filter_ready = pes_0_6_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_6_io_ifmap_ready = pes_0_6_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_6_io_pSum_ready = pes_0_6_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_8_clock = clock;
  assign NoC_0_8_reset = reset;
  assign NoC_0_8_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_8_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_8_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_8_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_8_io_dataPackageOut_ready = dss_0_7_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_7_clock = clock;
  assign pes_0_7_reset = reset;
  assign pes_0_7_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_7_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_7_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_7_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_7_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_7_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_7_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_7_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_7_io_filter_valid = dss_0_7_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_7_io_filter_bits = dss_0_7_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_7_io_ifmap_valid = dss_0_7_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_7_io_ifmap_bits = dss_0_7_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_7_io_pSumIn_valid = dss_0_7_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_7_io_pSumIn_bits = {{4{dss_0_7_io_pSum_bits[15]}},dss_0_7_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_7_io_pSumOut_ready = pes_1_7_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_7_io_dataIn_valid = NoC_0_8_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_7_io_dataIn_bits_data = {{11{NoC_0_8_io_dataPackageOut_bits_data[4]}},NoC_0_8_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_0_7_io_dataIn_bits_dataType = NoC_0_8_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_7_io_filter_ready = pes_0_7_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_7_io_ifmap_ready = pes_0_7_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_7_io_pSum_ready = pes_0_7_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_9_clock = clock;
  assign NoC_0_9_reset = reset;
  assign NoC_0_9_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_9_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_9_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_9_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_9_io_dataPackageOut_ready = dss_0_8_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_8_clock = clock;
  assign pes_0_8_reset = reset;
  assign pes_0_8_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_8_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_8_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_8_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_8_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_8_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_8_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_8_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_8_io_filter_valid = dss_0_8_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_8_io_filter_bits = dss_0_8_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_8_io_ifmap_valid = dss_0_8_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_8_io_ifmap_bits = dss_0_8_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_8_io_pSumIn_valid = dss_0_8_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_8_io_pSumIn_bits = {{4{dss_0_8_io_pSum_bits[15]}},dss_0_8_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_8_io_pSumOut_ready = pes_1_8_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_8_io_dataIn_valid = NoC_0_9_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_8_io_dataIn_bits_data = {{11{NoC_0_9_io_dataPackageOut_bits_data[4]}},NoC_0_9_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_0_8_io_dataIn_bits_dataType = NoC_0_9_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_8_io_filter_ready = pes_0_8_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_8_io_ifmap_ready = pes_0_8_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_8_io_pSum_ready = pes_0_8_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_10_clock = clock;
  assign NoC_0_10_reset = reset;
  assign NoC_0_10_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_10_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_10_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_10_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_10_io_dataPackageOut_ready = dss_0_9_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_9_clock = clock;
  assign pes_0_9_reset = reset;
  assign pes_0_9_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_9_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_9_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_9_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_9_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_9_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_9_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_9_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_9_io_filter_valid = dss_0_9_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_9_io_filter_bits = dss_0_9_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_9_io_ifmap_valid = dss_0_9_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_9_io_ifmap_bits = dss_0_9_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_9_io_pSumIn_valid = dss_0_9_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_9_io_pSumIn_bits = {{4{dss_0_9_io_pSum_bits[15]}},dss_0_9_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_9_io_pSumOut_ready = pes_1_9_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_9_io_dataIn_valid = NoC_0_10_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_9_io_dataIn_bits_data = {{11{NoC_0_10_io_dataPackageOut_bits_data[4]}},
    NoC_0_10_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_9_io_dataIn_bits_dataType = NoC_0_10_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_9_io_filter_ready = pes_0_9_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_9_io_ifmap_ready = pes_0_9_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_9_io_pSum_ready = pes_0_9_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_11_clock = clock;
  assign NoC_0_11_reset = reset;
  assign NoC_0_11_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_11_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_11_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_11_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_11_io_dataPackageOut_ready = dss_0_10_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_10_clock = clock;
  assign pes_0_10_reset = reset;
  assign pes_0_10_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_10_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_10_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_10_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_10_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_10_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_10_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_10_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_10_io_filter_valid = dss_0_10_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_10_io_filter_bits = dss_0_10_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_10_io_ifmap_valid = dss_0_10_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_10_io_ifmap_bits = dss_0_10_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_10_io_pSumIn_valid = dss_0_10_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_10_io_pSumIn_bits = {{4{dss_0_10_io_pSum_bits[15]}},dss_0_10_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_10_io_pSumOut_ready = pes_1_10_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_10_io_dataIn_valid = NoC_0_11_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_10_io_dataIn_bits_data = {{11{NoC_0_11_io_dataPackageOut_bits_data[4]}},
    NoC_0_11_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_10_io_dataIn_bits_dataType = NoC_0_11_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_10_io_filter_ready = pes_0_10_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_10_io_ifmap_ready = pes_0_10_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_10_io_pSum_ready = pes_0_10_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_12_clock = clock;
  assign NoC_0_12_reset = reset;
  assign NoC_0_12_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_12_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_12_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_12_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_12_io_dataPackageOut_ready = dss_0_11_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_11_clock = clock;
  assign pes_0_11_reset = reset;
  assign pes_0_11_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_11_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_11_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_11_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_11_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_11_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_11_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_11_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_11_io_filter_valid = dss_0_11_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_11_io_filter_bits = dss_0_11_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_11_io_ifmap_valid = dss_0_11_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_11_io_ifmap_bits = dss_0_11_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_11_io_pSumIn_valid = dss_0_11_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_11_io_pSumIn_bits = {{4{dss_0_11_io_pSum_bits[15]}},dss_0_11_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_11_io_pSumOut_ready = pes_1_11_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_11_io_dataIn_valid = NoC_0_12_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_11_io_dataIn_bits_data = {{11{NoC_0_12_io_dataPackageOut_bits_data[4]}},
    NoC_0_12_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_11_io_dataIn_bits_dataType = NoC_0_12_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_11_io_filter_ready = pes_0_11_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_11_io_ifmap_ready = pes_0_11_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_11_io_pSum_ready = pes_0_11_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_13_clock = clock;
  assign NoC_0_13_reset = reset;
  assign NoC_0_13_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_13_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_13_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_13_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_13_io_dataPackageOut_ready = dss_0_12_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_12_clock = clock;
  assign pes_0_12_reset = reset;
  assign pes_0_12_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_12_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_12_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_12_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_12_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_12_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_12_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_12_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_12_io_filter_valid = dss_0_12_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_12_io_filter_bits = dss_0_12_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_12_io_ifmap_valid = dss_0_12_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_12_io_ifmap_bits = dss_0_12_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_12_io_pSumIn_valid = dss_0_12_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_12_io_pSumIn_bits = {{4{dss_0_12_io_pSum_bits[15]}},dss_0_12_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_12_io_pSumOut_ready = pes_1_12_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_12_io_dataIn_valid = NoC_0_13_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_12_io_dataIn_bits_data = {{11{NoC_0_13_io_dataPackageOut_bits_data[4]}},
    NoC_0_13_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_12_io_dataIn_bits_dataType = NoC_0_13_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_12_io_filter_ready = pes_0_12_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_12_io_ifmap_ready = pes_0_12_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_12_io_pSum_ready = pes_0_12_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_14_clock = clock;
  assign NoC_0_14_reset = reset;
  assign NoC_0_14_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_14_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_14_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_14_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_14_io_dataPackageOut_ready = dss_0_13_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_13_clock = clock;
  assign pes_0_13_reset = reset;
  assign pes_0_13_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_13_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_13_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_13_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_13_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_13_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_13_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_13_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_13_io_filter_valid = dss_0_13_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_13_io_filter_bits = dss_0_13_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_13_io_ifmap_valid = dss_0_13_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_13_io_ifmap_bits = dss_0_13_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_13_io_pSumIn_valid = dss_0_13_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_13_io_pSumIn_bits = {{4{dss_0_13_io_pSum_bits[15]}},dss_0_13_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_13_io_pSumOut_ready = pes_1_13_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_13_io_dataIn_valid = NoC_0_14_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_13_io_dataIn_bits_data = {{11{NoC_0_14_io_dataPackageOut_bits_data[4]}},
    NoC_0_14_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_13_io_dataIn_bits_dataType = NoC_0_14_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_13_io_filter_ready = pes_0_13_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_13_io_ifmap_ready = pes_0_13_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_13_io_pSum_ready = pes_0_13_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_15_clock = clock;
  assign NoC_0_15_reset = reset;
  assign NoC_0_15_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_15_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_15_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_15_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_15_io_dataPackageOut_ready = dss_0_14_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_14_clock = clock;
  assign pes_0_14_reset = reset;
  assign pes_0_14_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_14_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_14_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_14_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_14_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_14_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_14_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_14_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_14_io_filter_valid = dss_0_14_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_14_io_filter_bits = dss_0_14_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_14_io_ifmap_valid = dss_0_14_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_14_io_ifmap_bits = dss_0_14_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_14_io_pSumIn_valid = dss_0_14_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_14_io_pSumIn_bits = {{4{dss_0_14_io_pSum_bits[15]}},dss_0_14_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_14_io_pSumOut_ready = pes_1_14_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_14_io_dataIn_valid = NoC_0_15_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_14_io_dataIn_bits_data = {{11{NoC_0_15_io_dataPackageOut_bits_data[4]}},
    NoC_0_15_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_14_io_dataIn_bits_dataType = NoC_0_15_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_14_io_filter_ready = pes_0_14_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_14_io_ifmap_ready = pes_0_14_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_14_io_pSum_ready = pes_0_14_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_16_clock = clock;
  assign NoC_0_16_reset = reset;
  assign NoC_0_16_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_16_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_16_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_16_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_16_io_dataPackageOut_ready = dss_0_15_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_15_clock = clock;
  assign pes_0_15_reset = reset;
  assign pes_0_15_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_15_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_15_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_15_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_15_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_15_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_15_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_15_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_15_io_filter_valid = dss_0_15_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_15_io_filter_bits = dss_0_15_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_15_io_ifmap_valid = dss_0_15_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_15_io_ifmap_bits = dss_0_15_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_15_io_pSumIn_valid = dss_0_15_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_15_io_pSumIn_bits = {{4{dss_0_15_io_pSum_bits[15]}},dss_0_15_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_15_io_pSumOut_ready = pes_1_15_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_15_io_dataIn_valid = NoC_0_16_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_15_io_dataIn_bits_data = {{11{NoC_0_16_io_dataPackageOut_bits_data[4]}},
    NoC_0_16_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_15_io_dataIn_bits_dataType = NoC_0_16_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_15_io_filter_ready = pes_0_15_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_15_io_ifmap_ready = pes_0_15_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_15_io_pSum_ready = pes_0_15_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_17_clock = clock;
  assign NoC_0_17_reset = reset;
  assign NoC_0_17_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_17_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_17_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_17_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_17_io_dataPackageOut_ready = dss_0_16_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_16_clock = clock;
  assign pes_0_16_reset = reset;
  assign pes_0_16_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_16_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_16_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_16_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_16_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_16_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_16_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_16_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_16_io_filter_valid = dss_0_16_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_16_io_filter_bits = dss_0_16_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_16_io_ifmap_valid = dss_0_16_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_16_io_ifmap_bits = dss_0_16_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_16_io_pSumIn_valid = dss_0_16_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_16_io_pSumIn_bits = {{4{dss_0_16_io_pSum_bits[15]}},dss_0_16_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_16_io_pSumOut_ready = pes_1_16_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_16_io_dataIn_valid = NoC_0_17_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_16_io_dataIn_bits_data = {{11{NoC_0_17_io_dataPackageOut_bits_data[4]}},
    NoC_0_17_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_16_io_dataIn_bits_dataType = NoC_0_17_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_16_io_filter_ready = pes_0_16_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_16_io_ifmap_ready = pes_0_16_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_16_io_pSum_ready = pes_0_16_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_18_clock = clock;
  assign NoC_0_18_reset = reset;
  assign NoC_0_18_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_18_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_18_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_18_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_18_io_dataPackageOut_ready = dss_0_17_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_17_clock = clock;
  assign pes_0_17_reset = reset;
  assign pes_0_17_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_17_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_17_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_17_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_17_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_17_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_17_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_17_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_17_io_filter_valid = dss_0_17_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_17_io_filter_bits = dss_0_17_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_17_io_ifmap_valid = dss_0_17_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_17_io_ifmap_bits = dss_0_17_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_17_io_pSumIn_valid = dss_0_17_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_17_io_pSumIn_bits = {{4{dss_0_17_io_pSum_bits[15]}},dss_0_17_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_17_io_pSumOut_ready = pes_1_17_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_17_io_dataIn_valid = NoC_0_18_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_17_io_dataIn_bits_data = {{11{NoC_0_18_io_dataPackageOut_bits_data[4]}},
    NoC_0_18_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_17_io_dataIn_bits_dataType = NoC_0_18_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_17_io_filter_ready = pes_0_17_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_17_io_ifmap_ready = pes_0_17_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_17_io_pSum_ready = pes_0_17_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_19_clock = clock;
  assign NoC_0_19_reset = reset;
  assign NoC_0_19_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_19_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_19_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_19_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_19_io_dataPackageOut_ready = dss_0_18_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_18_clock = clock;
  assign pes_0_18_reset = reset;
  assign pes_0_18_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_18_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_18_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_18_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_18_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_18_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_18_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_18_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_18_io_filter_valid = dss_0_18_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_18_io_filter_bits = dss_0_18_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_18_io_ifmap_valid = dss_0_18_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_18_io_ifmap_bits = dss_0_18_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_18_io_pSumIn_valid = dss_0_18_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_18_io_pSumIn_bits = {{4{dss_0_18_io_pSum_bits[15]}},dss_0_18_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_18_io_pSumOut_ready = pes_1_18_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_18_io_dataIn_valid = NoC_0_19_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_18_io_dataIn_bits_data = {{11{NoC_0_19_io_dataPackageOut_bits_data[4]}},
    NoC_0_19_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_18_io_dataIn_bits_dataType = NoC_0_19_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_18_io_filter_ready = pes_0_18_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_18_io_ifmap_ready = pes_0_18_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_18_io_pSum_ready = pes_0_18_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_20_clock = clock;
  assign NoC_0_20_reset = reset;
  assign NoC_0_20_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_20_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_20_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_20_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_20_io_dataPackageOut_ready = dss_0_19_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_19_clock = clock;
  assign pes_0_19_reset = reset;
  assign pes_0_19_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_19_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_19_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_19_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_19_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_19_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_19_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_19_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_19_io_filter_valid = dss_0_19_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_19_io_filter_bits = dss_0_19_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_19_io_ifmap_valid = dss_0_19_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_19_io_ifmap_bits = dss_0_19_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_19_io_pSumIn_valid = dss_0_19_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_19_io_pSumIn_bits = {{4{dss_0_19_io_pSum_bits[15]}},dss_0_19_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_19_io_pSumOut_ready = pes_1_19_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_19_io_dataIn_valid = NoC_0_20_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_19_io_dataIn_bits_data = {{11{NoC_0_20_io_dataPackageOut_bits_data[4]}},
    NoC_0_20_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_19_io_dataIn_bits_dataType = NoC_0_20_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_19_io_filter_ready = pes_0_19_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_19_io_ifmap_ready = pes_0_19_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_19_io_pSum_ready = pes_0_19_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_21_clock = clock;
  assign NoC_0_21_reset = reset;
  assign NoC_0_21_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_21_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_21_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_21_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_21_io_dataPackageOut_ready = dss_0_20_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_20_clock = clock;
  assign pes_0_20_reset = reset;
  assign pes_0_20_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_20_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_20_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_20_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_20_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_20_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_20_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_20_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_20_io_filter_valid = dss_0_20_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_20_io_filter_bits = dss_0_20_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_20_io_ifmap_valid = dss_0_20_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_20_io_ifmap_bits = dss_0_20_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_20_io_pSumIn_valid = dss_0_20_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_20_io_pSumIn_bits = {{4{dss_0_20_io_pSum_bits[15]}},dss_0_20_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_20_io_pSumOut_ready = pes_1_20_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_20_io_dataIn_valid = NoC_0_21_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_20_io_dataIn_bits_data = {{11{NoC_0_21_io_dataPackageOut_bits_data[4]}},
    NoC_0_21_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_20_io_dataIn_bits_dataType = NoC_0_21_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_20_io_filter_ready = pes_0_20_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_20_io_ifmap_ready = pes_0_20_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_20_io_pSum_ready = pes_0_20_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_22_clock = clock;
  assign NoC_0_22_reset = reset;
  assign NoC_0_22_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_22_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_22_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_22_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_22_io_dataPackageOut_ready = dss_0_21_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_21_clock = clock;
  assign pes_0_21_reset = reset;
  assign pes_0_21_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_21_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_21_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_21_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_21_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_21_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_21_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_21_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_21_io_filter_valid = dss_0_21_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_21_io_filter_bits = dss_0_21_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_21_io_ifmap_valid = dss_0_21_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_21_io_ifmap_bits = dss_0_21_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_21_io_pSumIn_valid = dss_0_21_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_21_io_pSumIn_bits = {{4{dss_0_21_io_pSum_bits[15]}},dss_0_21_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_21_io_pSumOut_ready = pes_1_21_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_21_io_dataIn_valid = NoC_0_22_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_21_io_dataIn_bits_data = {{11{NoC_0_22_io_dataPackageOut_bits_data[4]}},
    NoC_0_22_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_21_io_dataIn_bits_dataType = NoC_0_22_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_21_io_filter_ready = pes_0_21_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_21_io_ifmap_ready = pes_0_21_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_21_io_pSum_ready = pes_0_21_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_23_clock = clock;
  assign NoC_0_23_reset = reset;
  assign NoC_0_23_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_23_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_23_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_23_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_23_io_dataPackageOut_ready = dss_0_22_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_22_clock = clock;
  assign pes_0_22_reset = reset;
  assign pes_0_22_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_22_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_22_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_22_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_22_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_22_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_22_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_22_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_22_io_filter_valid = dss_0_22_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_22_io_filter_bits = dss_0_22_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_22_io_ifmap_valid = dss_0_22_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_22_io_ifmap_bits = dss_0_22_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_22_io_pSumIn_valid = dss_0_22_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_22_io_pSumIn_bits = {{4{dss_0_22_io_pSum_bits[15]}},dss_0_22_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_22_io_pSumOut_ready = pes_1_22_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_22_io_dataIn_valid = NoC_0_23_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_22_io_dataIn_bits_data = {{11{NoC_0_23_io_dataPackageOut_bits_data[4]}},
    NoC_0_23_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_22_io_dataIn_bits_dataType = NoC_0_23_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_22_io_filter_ready = pes_0_22_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_22_io_ifmap_ready = pes_0_22_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_22_io_pSum_ready = pes_0_22_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_0_24_clock = clock;
  assign NoC_0_24_reset = reset;
  assign NoC_0_24_io_dataPackageIn_valid = NoC_0_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_0_24_io_dataPackageIn_bits_data = NoC_0_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_0_24_io_dataPackageIn_bits_dataType = NoC_0_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_0_24_io_dataPackageIn_bits_positon_col = NoC_0_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_0_24_io_dataPackageOut_ready = dss_0_23_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_0_23_clock = clock;
  assign pes_0_23_reset = reset;
  assign pes_0_23_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_0_23_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_0_23_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_0_23_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_0_23_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_0_23_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_0_23_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_0_23_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_0_23_io_filter_valid = dss_0_23_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_0_23_io_filter_bits = dss_0_23_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_0_23_io_ifmap_valid = dss_0_23_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_0_23_io_ifmap_bits = dss_0_23_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_0_23_io_pSumIn_valid = dss_0_23_io_pSum_valid; // @[PEArray.scala 46:24]
  assign pes_0_23_io_pSumIn_bits = {{4{dss_0_23_io_pSum_bits[15]}},dss_0_23_io_pSum_bits}; // @[PEArray.scala 46:24]
  assign pes_0_23_io_pSumOut_ready = pes_1_23_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_0_23_io_dataIn_valid = NoC_0_24_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_0_23_io_dataIn_bits_data = {{11{NoC_0_24_io_dataPackageOut_bits_data[4]}},
    NoC_0_24_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_0_23_io_dataIn_bits_dataType = NoC_0_24_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_0_23_io_filter_ready = pes_0_23_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_0_23_io_ifmap_ready = pes_0_23_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_0_23_io_pSum_ready = pes_0_23_io_pSumIn_ready; // @[PEArray.scala 46:24]
  assign NoC_1_0_clock = clock;
  assign NoC_1_0_reset = reset;
  assign NoC_1_0_io_dataPackageIn_valid = io_dataIn_valid; // @[PEArray.scala 84:35]
  assign NoC_1_0_io_dataPackageIn_bits_data = io_dataIn_bits_data; // @[PEArray.scala 85:34]
  assign NoC_1_0_io_dataPackageIn_bits_dataType = io_dataIn_bits_dataType; // @[PEArray.scala 85:34]
  assign NoC_1_0_io_dataPackageIn_bits_positon_row = io_dataIn_bits_positon_row; // @[PEArray.scala 85:34]
  assign NoC_1_0_io_dataPackageIn_bits_positon_col = io_dataIn_bits_positon_col; // @[PEArray.scala 85:34]
  assign NoC_1_0_io_dataPackageOut_ready = NoC_1_1_io_dataPackageIn_ready | NoC_1_2_io_dataPackageIn_ready |
    NoC_1_3_io_dataPackageIn_ready | NoC_1_4_io_dataPackageIn_ready | NoC_1_5_io_dataPackageIn_ready |
    NoC_1_6_io_dataPackageIn_ready | NoC_1_7_io_dataPackageIn_ready | NoC_1_8_io_dataPackageIn_ready |
    NoC_1_9_io_dataPackageIn_ready | NoC_1_10_io_dataPackageIn_ready | NoC_1_11_io_dataPackageIn_ready |
    NoC_1_12_io_dataPackageIn_ready | NoC_1_13_io_dataPackageIn_ready | NoC_1_14_io_dataPackageIn_ready |
    NoC_1_15_io_dataPackageIn_ready | NoC_1_16_io_dataPackageIn_ready | NoC_1_17_io_dataPackageIn_ready |
    NoC_1_18_io_dataPackageIn_ready | NoC_1_19_io_dataPackageIn_ready | NoC_1_20_io_dataPackageIn_ready |
    NoC_1_21_io_dataPackageIn_ready | NoC_1_22_io_dataPackageIn_ready | NoC_1_23_io_dataPackageIn_ready |
    NoC_1_24_io_dataPackageIn_ready; // @[PEArray.scala 83:17]
  assign NoC_1_1_clock = clock;
  assign NoC_1_1_reset = reset;
  assign NoC_1_1_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_1_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_1_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_1_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_1_io_dataPackageOut_ready = dss_1_0_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_0_clock = clock;
  assign pes_1_0_reset = reset;
  assign pes_1_0_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_0_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_0_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_0_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_0_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_0_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_0_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_0_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_0_io_filter_valid = dss_1_0_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_0_io_filter_bits = dss_1_0_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_0_io_ifmap_valid = dss_1_0_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_0_io_ifmap_bits = dss_1_0_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_0_io_pSumIn_valid = pes_0_0_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_0_io_pSumIn_bits = pes_0_0_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_0_io_pSumOut_ready = pes_2_0_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_0_io_dataIn_valid = NoC_1_1_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_0_io_dataIn_bits_data = {{11{NoC_1_1_io_dataPackageOut_bits_data[4]}},NoC_1_1_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_1_0_io_dataIn_bits_dataType = NoC_1_1_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_0_io_filter_ready = pes_1_0_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_0_io_ifmap_ready = pes_1_0_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_0_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_2_clock = clock;
  assign NoC_1_2_reset = reset;
  assign NoC_1_2_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_2_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_2_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_2_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_2_io_dataPackageOut_ready = dss_1_1_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_1_clock = clock;
  assign pes_1_1_reset = reset;
  assign pes_1_1_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_1_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_1_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_1_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_1_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_1_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_1_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_1_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_1_io_filter_valid = dss_1_1_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_1_io_filter_bits = dss_1_1_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_1_io_ifmap_valid = dss_1_1_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_1_io_ifmap_bits = dss_1_1_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_1_io_pSumIn_valid = pes_0_1_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_1_io_pSumIn_bits = pes_0_1_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_1_io_pSumOut_ready = pes_2_1_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_1_io_dataIn_valid = NoC_1_2_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_1_io_dataIn_bits_data = {{11{NoC_1_2_io_dataPackageOut_bits_data[4]}},NoC_1_2_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_1_1_io_dataIn_bits_dataType = NoC_1_2_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_1_io_filter_ready = pes_1_1_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_1_io_ifmap_ready = pes_1_1_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_1_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_3_clock = clock;
  assign NoC_1_3_reset = reset;
  assign NoC_1_3_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_3_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_3_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_3_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_3_io_dataPackageOut_ready = dss_1_2_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_2_clock = clock;
  assign pes_1_2_reset = reset;
  assign pes_1_2_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_2_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_2_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_2_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_2_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_2_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_2_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_2_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_2_io_filter_valid = dss_1_2_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_2_io_filter_bits = dss_1_2_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_2_io_ifmap_valid = dss_1_2_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_2_io_ifmap_bits = dss_1_2_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_2_io_pSumIn_valid = pes_0_2_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_2_io_pSumIn_bits = pes_0_2_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_2_io_pSumOut_ready = pes_2_2_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_2_io_dataIn_valid = NoC_1_3_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_2_io_dataIn_bits_data = {{11{NoC_1_3_io_dataPackageOut_bits_data[4]}},NoC_1_3_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_1_2_io_dataIn_bits_dataType = NoC_1_3_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_2_io_filter_ready = pes_1_2_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_2_io_ifmap_ready = pes_1_2_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_2_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_4_clock = clock;
  assign NoC_1_4_reset = reset;
  assign NoC_1_4_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_4_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_4_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_4_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_4_io_dataPackageOut_ready = dss_1_3_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_3_clock = clock;
  assign pes_1_3_reset = reset;
  assign pes_1_3_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_3_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_3_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_3_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_3_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_3_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_3_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_3_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_3_io_filter_valid = dss_1_3_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_3_io_filter_bits = dss_1_3_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_3_io_ifmap_valid = dss_1_3_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_3_io_ifmap_bits = dss_1_3_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_3_io_pSumIn_valid = pes_0_3_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_3_io_pSumIn_bits = pes_0_3_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_3_io_pSumOut_ready = pes_2_3_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_3_io_dataIn_valid = NoC_1_4_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_3_io_dataIn_bits_data = {{11{NoC_1_4_io_dataPackageOut_bits_data[4]}},NoC_1_4_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_1_3_io_dataIn_bits_dataType = NoC_1_4_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_3_io_filter_ready = pes_1_3_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_3_io_ifmap_ready = pes_1_3_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_3_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_5_clock = clock;
  assign NoC_1_5_reset = reset;
  assign NoC_1_5_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_5_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_5_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_5_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_5_io_dataPackageOut_ready = dss_1_4_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_4_clock = clock;
  assign pes_1_4_reset = reset;
  assign pes_1_4_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_4_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_4_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_4_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_4_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_4_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_4_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_4_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_4_io_filter_valid = dss_1_4_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_4_io_filter_bits = dss_1_4_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_4_io_ifmap_valid = dss_1_4_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_4_io_ifmap_bits = dss_1_4_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_4_io_pSumIn_valid = pes_0_4_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_4_io_pSumIn_bits = pes_0_4_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_4_io_pSumOut_ready = pes_2_4_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_4_io_dataIn_valid = NoC_1_5_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_4_io_dataIn_bits_data = {{11{NoC_1_5_io_dataPackageOut_bits_data[4]}},NoC_1_5_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_1_4_io_dataIn_bits_dataType = NoC_1_5_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_4_io_filter_ready = pes_1_4_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_4_io_ifmap_ready = pes_1_4_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_4_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_6_clock = clock;
  assign NoC_1_6_reset = reset;
  assign NoC_1_6_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_6_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_6_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_6_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_6_io_dataPackageOut_ready = dss_1_5_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_5_clock = clock;
  assign pes_1_5_reset = reset;
  assign pes_1_5_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_5_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_5_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_5_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_5_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_5_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_5_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_5_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_5_io_filter_valid = dss_1_5_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_5_io_filter_bits = dss_1_5_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_5_io_ifmap_valid = dss_1_5_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_5_io_ifmap_bits = dss_1_5_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_5_io_pSumIn_valid = pes_0_5_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_5_io_pSumIn_bits = pes_0_5_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_5_io_pSumOut_ready = pes_2_5_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_5_io_dataIn_valid = NoC_1_6_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_5_io_dataIn_bits_data = {{11{NoC_1_6_io_dataPackageOut_bits_data[4]}},NoC_1_6_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_1_5_io_dataIn_bits_dataType = NoC_1_6_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_5_io_filter_ready = pes_1_5_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_5_io_ifmap_ready = pes_1_5_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_5_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_7_clock = clock;
  assign NoC_1_7_reset = reset;
  assign NoC_1_7_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_7_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_7_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_7_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_7_io_dataPackageOut_ready = dss_1_6_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_6_clock = clock;
  assign pes_1_6_reset = reset;
  assign pes_1_6_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_6_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_6_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_6_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_6_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_6_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_6_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_6_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_6_io_filter_valid = dss_1_6_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_6_io_filter_bits = dss_1_6_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_6_io_ifmap_valid = dss_1_6_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_6_io_ifmap_bits = dss_1_6_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_6_io_pSumIn_valid = pes_0_6_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_6_io_pSumIn_bits = pes_0_6_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_6_io_pSumOut_ready = pes_2_6_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_6_io_dataIn_valid = NoC_1_7_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_6_io_dataIn_bits_data = {{11{NoC_1_7_io_dataPackageOut_bits_data[4]}},NoC_1_7_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_1_6_io_dataIn_bits_dataType = NoC_1_7_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_6_io_filter_ready = pes_1_6_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_6_io_ifmap_ready = pes_1_6_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_6_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_8_clock = clock;
  assign NoC_1_8_reset = reset;
  assign NoC_1_8_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_8_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_8_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_8_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_8_io_dataPackageOut_ready = dss_1_7_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_7_clock = clock;
  assign pes_1_7_reset = reset;
  assign pes_1_7_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_7_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_7_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_7_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_7_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_7_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_7_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_7_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_7_io_filter_valid = dss_1_7_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_7_io_filter_bits = dss_1_7_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_7_io_ifmap_valid = dss_1_7_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_7_io_ifmap_bits = dss_1_7_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_7_io_pSumIn_valid = pes_0_7_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_7_io_pSumIn_bits = pes_0_7_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_7_io_pSumOut_ready = pes_2_7_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_7_io_dataIn_valid = NoC_1_8_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_7_io_dataIn_bits_data = {{11{NoC_1_8_io_dataPackageOut_bits_data[4]}},NoC_1_8_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_1_7_io_dataIn_bits_dataType = NoC_1_8_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_7_io_filter_ready = pes_1_7_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_7_io_ifmap_ready = pes_1_7_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_7_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_9_clock = clock;
  assign NoC_1_9_reset = reset;
  assign NoC_1_9_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_9_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_9_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_9_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_9_io_dataPackageOut_ready = dss_1_8_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_8_clock = clock;
  assign pes_1_8_reset = reset;
  assign pes_1_8_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_8_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_8_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_8_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_8_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_8_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_8_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_8_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_8_io_filter_valid = dss_1_8_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_8_io_filter_bits = dss_1_8_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_8_io_ifmap_valid = dss_1_8_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_8_io_ifmap_bits = dss_1_8_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_8_io_pSumIn_valid = pes_0_8_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_8_io_pSumIn_bits = pes_0_8_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_8_io_pSumOut_ready = pes_2_8_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_8_io_dataIn_valid = NoC_1_9_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_8_io_dataIn_bits_data = {{11{NoC_1_9_io_dataPackageOut_bits_data[4]}},NoC_1_9_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_1_8_io_dataIn_bits_dataType = NoC_1_9_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_8_io_filter_ready = pes_1_8_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_8_io_ifmap_ready = pes_1_8_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_8_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_10_clock = clock;
  assign NoC_1_10_reset = reset;
  assign NoC_1_10_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_10_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_10_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_10_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_10_io_dataPackageOut_ready = dss_1_9_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_9_clock = clock;
  assign pes_1_9_reset = reset;
  assign pes_1_9_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_9_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_9_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_9_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_9_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_9_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_9_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_9_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_9_io_filter_valid = dss_1_9_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_9_io_filter_bits = dss_1_9_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_9_io_ifmap_valid = dss_1_9_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_9_io_ifmap_bits = dss_1_9_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_9_io_pSumIn_valid = pes_0_9_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_9_io_pSumIn_bits = pes_0_9_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_9_io_pSumOut_ready = pes_2_9_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_9_io_dataIn_valid = NoC_1_10_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_9_io_dataIn_bits_data = {{11{NoC_1_10_io_dataPackageOut_bits_data[4]}},
    NoC_1_10_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_9_io_dataIn_bits_dataType = NoC_1_10_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_9_io_filter_ready = pes_1_9_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_9_io_ifmap_ready = pes_1_9_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_9_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_11_clock = clock;
  assign NoC_1_11_reset = reset;
  assign NoC_1_11_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_11_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_11_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_11_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_11_io_dataPackageOut_ready = dss_1_10_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_10_clock = clock;
  assign pes_1_10_reset = reset;
  assign pes_1_10_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_10_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_10_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_10_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_10_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_10_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_10_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_10_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_10_io_filter_valid = dss_1_10_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_10_io_filter_bits = dss_1_10_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_10_io_ifmap_valid = dss_1_10_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_10_io_ifmap_bits = dss_1_10_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_10_io_pSumIn_valid = pes_0_10_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_10_io_pSumIn_bits = pes_0_10_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_10_io_pSumOut_ready = pes_2_10_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_10_io_dataIn_valid = NoC_1_11_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_10_io_dataIn_bits_data = {{11{NoC_1_11_io_dataPackageOut_bits_data[4]}},
    NoC_1_11_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_10_io_dataIn_bits_dataType = NoC_1_11_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_10_io_filter_ready = pes_1_10_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_10_io_ifmap_ready = pes_1_10_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_10_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_12_clock = clock;
  assign NoC_1_12_reset = reset;
  assign NoC_1_12_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_12_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_12_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_12_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_12_io_dataPackageOut_ready = dss_1_11_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_11_clock = clock;
  assign pes_1_11_reset = reset;
  assign pes_1_11_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_11_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_11_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_11_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_11_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_11_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_11_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_11_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_11_io_filter_valid = dss_1_11_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_11_io_filter_bits = dss_1_11_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_11_io_ifmap_valid = dss_1_11_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_11_io_ifmap_bits = dss_1_11_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_11_io_pSumIn_valid = pes_0_11_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_11_io_pSumIn_bits = pes_0_11_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_11_io_pSumOut_ready = pes_2_11_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_11_io_dataIn_valid = NoC_1_12_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_11_io_dataIn_bits_data = {{11{NoC_1_12_io_dataPackageOut_bits_data[4]}},
    NoC_1_12_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_11_io_dataIn_bits_dataType = NoC_1_12_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_11_io_filter_ready = pes_1_11_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_11_io_ifmap_ready = pes_1_11_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_11_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_13_clock = clock;
  assign NoC_1_13_reset = reset;
  assign NoC_1_13_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_13_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_13_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_13_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_13_io_dataPackageOut_ready = dss_1_12_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_12_clock = clock;
  assign pes_1_12_reset = reset;
  assign pes_1_12_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_12_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_12_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_12_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_12_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_12_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_12_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_12_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_12_io_filter_valid = dss_1_12_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_12_io_filter_bits = dss_1_12_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_12_io_ifmap_valid = dss_1_12_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_12_io_ifmap_bits = dss_1_12_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_12_io_pSumIn_valid = pes_0_12_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_12_io_pSumIn_bits = pes_0_12_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_12_io_pSumOut_ready = pes_2_12_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_12_io_dataIn_valid = NoC_1_13_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_12_io_dataIn_bits_data = {{11{NoC_1_13_io_dataPackageOut_bits_data[4]}},
    NoC_1_13_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_12_io_dataIn_bits_dataType = NoC_1_13_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_12_io_filter_ready = pes_1_12_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_12_io_ifmap_ready = pes_1_12_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_12_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_14_clock = clock;
  assign NoC_1_14_reset = reset;
  assign NoC_1_14_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_14_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_14_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_14_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_14_io_dataPackageOut_ready = dss_1_13_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_13_clock = clock;
  assign pes_1_13_reset = reset;
  assign pes_1_13_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_13_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_13_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_13_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_13_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_13_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_13_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_13_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_13_io_filter_valid = dss_1_13_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_13_io_filter_bits = dss_1_13_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_13_io_ifmap_valid = dss_1_13_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_13_io_ifmap_bits = dss_1_13_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_13_io_pSumIn_valid = pes_0_13_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_13_io_pSumIn_bits = pes_0_13_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_13_io_pSumOut_ready = pes_2_13_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_13_io_dataIn_valid = NoC_1_14_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_13_io_dataIn_bits_data = {{11{NoC_1_14_io_dataPackageOut_bits_data[4]}},
    NoC_1_14_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_13_io_dataIn_bits_dataType = NoC_1_14_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_13_io_filter_ready = pes_1_13_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_13_io_ifmap_ready = pes_1_13_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_13_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_15_clock = clock;
  assign NoC_1_15_reset = reset;
  assign NoC_1_15_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_15_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_15_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_15_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_15_io_dataPackageOut_ready = dss_1_14_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_14_clock = clock;
  assign pes_1_14_reset = reset;
  assign pes_1_14_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_14_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_14_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_14_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_14_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_14_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_14_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_14_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_14_io_filter_valid = dss_1_14_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_14_io_filter_bits = dss_1_14_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_14_io_ifmap_valid = dss_1_14_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_14_io_ifmap_bits = dss_1_14_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_14_io_pSumIn_valid = pes_0_14_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_14_io_pSumIn_bits = pes_0_14_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_14_io_pSumOut_ready = pes_2_14_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_14_io_dataIn_valid = NoC_1_15_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_14_io_dataIn_bits_data = {{11{NoC_1_15_io_dataPackageOut_bits_data[4]}},
    NoC_1_15_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_14_io_dataIn_bits_dataType = NoC_1_15_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_14_io_filter_ready = pes_1_14_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_14_io_ifmap_ready = pes_1_14_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_14_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_16_clock = clock;
  assign NoC_1_16_reset = reset;
  assign NoC_1_16_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_16_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_16_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_16_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_16_io_dataPackageOut_ready = dss_1_15_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_15_clock = clock;
  assign pes_1_15_reset = reset;
  assign pes_1_15_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_15_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_15_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_15_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_15_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_15_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_15_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_15_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_15_io_filter_valid = dss_1_15_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_15_io_filter_bits = dss_1_15_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_15_io_ifmap_valid = dss_1_15_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_15_io_ifmap_bits = dss_1_15_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_15_io_pSumIn_valid = pes_0_15_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_15_io_pSumIn_bits = pes_0_15_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_15_io_pSumOut_ready = pes_2_15_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_15_io_dataIn_valid = NoC_1_16_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_15_io_dataIn_bits_data = {{11{NoC_1_16_io_dataPackageOut_bits_data[4]}},
    NoC_1_16_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_15_io_dataIn_bits_dataType = NoC_1_16_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_15_io_filter_ready = pes_1_15_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_15_io_ifmap_ready = pes_1_15_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_15_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_17_clock = clock;
  assign NoC_1_17_reset = reset;
  assign NoC_1_17_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_17_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_17_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_17_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_17_io_dataPackageOut_ready = dss_1_16_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_16_clock = clock;
  assign pes_1_16_reset = reset;
  assign pes_1_16_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_16_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_16_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_16_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_16_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_16_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_16_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_16_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_16_io_filter_valid = dss_1_16_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_16_io_filter_bits = dss_1_16_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_16_io_ifmap_valid = dss_1_16_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_16_io_ifmap_bits = dss_1_16_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_16_io_pSumIn_valid = pes_0_16_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_16_io_pSumIn_bits = pes_0_16_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_16_io_pSumOut_ready = pes_2_16_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_16_io_dataIn_valid = NoC_1_17_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_16_io_dataIn_bits_data = {{11{NoC_1_17_io_dataPackageOut_bits_data[4]}},
    NoC_1_17_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_16_io_dataIn_bits_dataType = NoC_1_17_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_16_io_filter_ready = pes_1_16_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_16_io_ifmap_ready = pes_1_16_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_16_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_18_clock = clock;
  assign NoC_1_18_reset = reset;
  assign NoC_1_18_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_18_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_18_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_18_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_18_io_dataPackageOut_ready = dss_1_17_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_17_clock = clock;
  assign pes_1_17_reset = reset;
  assign pes_1_17_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_17_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_17_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_17_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_17_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_17_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_17_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_17_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_17_io_filter_valid = dss_1_17_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_17_io_filter_bits = dss_1_17_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_17_io_ifmap_valid = dss_1_17_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_17_io_ifmap_bits = dss_1_17_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_17_io_pSumIn_valid = pes_0_17_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_17_io_pSumIn_bits = pes_0_17_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_17_io_pSumOut_ready = pes_2_17_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_17_io_dataIn_valid = NoC_1_18_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_17_io_dataIn_bits_data = {{11{NoC_1_18_io_dataPackageOut_bits_data[4]}},
    NoC_1_18_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_17_io_dataIn_bits_dataType = NoC_1_18_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_17_io_filter_ready = pes_1_17_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_17_io_ifmap_ready = pes_1_17_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_17_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_19_clock = clock;
  assign NoC_1_19_reset = reset;
  assign NoC_1_19_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_19_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_19_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_19_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_19_io_dataPackageOut_ready = dss_1_18_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_18_clock = clock;
  assign pes_1_18_reset = reset;
  assign pes_1_18_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_18_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_18_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_18_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_18_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_18_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_18_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_18_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_18_io_filter_valid = dss_1_18_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_18_io_filter_bits = dss_1_18_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_18_io_ifmap_valid = dss_1_18_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_18_io_ifmap_bits = dss_1_18_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_18_io_pSumIn_valid = pes_0_18_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_18_io_pSumIn_bits = pes_0_18_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_18_io_pSumOut_ready = pes_2_18_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_18_io_dataIn_valid = NoC_1_19_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_18_io_dataIn_bits_data = {{11{NoC_1_19_io_dataPackageOut_bits_data[4]}},
    NoC_1_19_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_18_io_dataIn_bits_dataType = NoC_1_19_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_18_io_filter_ready = pes_1_18_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_18_io_ifmap_ready = pes_1_18_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_18_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_20_clock = clock;
  assign NoC_1_20_reset = reset;
  assign NoC_1_20_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_20_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_20_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_20_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_20_io_dataPackageOut_ready = dss_1_19_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_19_clock = clock;
  assign pes_1_19_reset = reset;
  assign pes_1_19_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_19_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_19_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_19_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_19_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_19_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_19_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_19_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_19_io_filter_valid = dss_1_19_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_19_io_filter_bits = dss_1_19_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_19_io_ifmap_valid = dss_1_19_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_19_io_ifmap_bits = dss_1_19_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_19_io_pSumIn_valid = pes_0_19_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_19_io_pSumIn_bits = pes_0_19_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_19_io_pSumOut_ready = pes_2_19_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_19_io_dataIn_valid = NoC_1_20_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_19_io_dataIn_bits_data = {{11{NoC_1_20_io_dataPackageOut_bits_data[4]}},
    NoC_1_20_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_19_io_dataIn_bits_dataType = NoC_1_20_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_19_io_filter_ready = pes_1_19_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_19_io_ifmap_ready = pes_1_19_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_19_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_21_clock = clock;
  assign NoC_1_21_reset = reset;
  assign NoC_1_21_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_21_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_21_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_21_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_21_io_dataPackageOut_ready = dss_1_20_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_20_clock = clock;
  assign pes_1_20_reset = reset;
  assign pes_1_20_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_20_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_20_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_20_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_20_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_20_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_20_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_20_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_20_io_filter_valid = dss_1_20_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_20_io_filter_bits = dss_1_20_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_20_io_ifmap_valid = dss_1_20_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_20_io_ifmap_bits = dss_1_20_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_20_io_pSumIn_valid = pes_0_20_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_20_io_pSumIn_bits = pes_0_20_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_20_io_pSumOut_ready = pes_2_20_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_20_io_dataIn_valid = NoC_1_21_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_20_io_dataIn_bits_data = {{11{NoC_1_21_io_dataPackageOut_bits_data[4]}},
    NoC_1_21_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_20_io_dataIn_bits_dataType = NoC_1_21_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_20_io_filter_ready = pes_1_20_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_20_io_ifmap_ready = pes_1_20_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_20_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_22_clock = clock;
  assign NoC_1_22_reset = reset;
  assign NoC_1_22_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_22_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_22_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_22_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_22_io_dataPackageOut_ready = dss_1_21_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_21_clock = clock;
  assign pes_1_21_reset = reset;
  assign pes_1_21_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_21_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_21_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_21_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_21_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_21_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_21_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_21_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_21_io_filter_valid = dss_1_21_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_21_io_filter_bits = dss_1_21_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_21_io_ifmap_valid = dss_1_21_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_21_io_ifmap_bits = dss_1_21_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_21_io_pSumIn_valid = pes_0_21_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_21_io_pSumIn_bits = pes_0_21_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_21_io_pSumOut_ready = pes_2_21_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_21_io_dataIn_valid = NoC_1_22_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_21_io_dataIn_bits_data = {{11{NoC_1_22_io_dataPackageOut_bits_data[4]}},
    NoC_1_22_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_21_io_dataIn_bits_dataType = NoC_1_22_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_21_io_filter_ready = pes_1_21_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_21_io_ifmap_ready = pes_1_21_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_21_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_23_clock = clock;
  assign NoC_1_23_reset = reset;
  assign NoC_1_23_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_23_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_23_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_23_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_23_io_dataPackageOut_ready = dss_1_22_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_22_clock = clock;
  assign pes_1_22_reset = reset;
  assign pes_1_22_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_22_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_22_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_22_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_22_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_22_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_22_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_22_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_22_io_filter_valid = dss_1_22_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_22_io_filter_bits = dss_1_22_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_22_io_ifmap_valid = dss_1_22_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_22_io_ifmap_bits = dss_1_22_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_22_io_pSumIn_valid = pes_0_22_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_22_io_pSumIn_bits = pes_0_22_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_22_io_pSumOut_ready = pes_2_22_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_22_io_dataIn_valid = NoC_1_23_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_22_io_dataIn_bits_data = {{11{NoC_1_23_io_dataPackageOut_bits_data[4]}},
    NoC_1_23_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_22_io_dataIn_bits_dataType = NoC_1_23_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_22_io_filter_ready = pes_1_22_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_22_io_ifmap_ready = pes_1_22_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_22_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_1_24_clock = clock;
  assign NoC_1_24_reset = reset;
  assign NoC_1_24_io_dataPackageIn_valid = NoC_1_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_1_24_io_dataPackageIn_bits_data = NoC_1_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_1_24_io_dataPackageIn_bits_dataType = NoC_1_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_1_24_io_dataPackageIn_bits_positon_col = NoC_1_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_1_24_io_dataPackageOut_ready = dss_1_23_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_1_23_clock = clock;
  assign pes_1_23_reset = reset;
  assign pes_1_23_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_1_23_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_1_23_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_1_23_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_1_23_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_1_23_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_1_23_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_1_23_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_1_23_io_filter_valid = dss_1_23_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_1_23_io_filter_bits = dss_1_23_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_1_23_io_ifmap_valid = dss_1_23_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_1_23_io_ifmap_bits = dss_1_23_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_1_23_io_pSumIn_valid = pes_0_23_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_1_23_io_pSumIn_bits = pes_0_23_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_1_23_io_pSumOut_ready = pes_2_23_io_pSumIn_ready; // @[PEArray.scala 93:27]
  assign dss_1_23_io_dataIn_valid = NoC_1_24_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_1_23_io_dataIn_bits_data = {{11{NoC_1_24_io_dataPackageOut_bits_data[4]}},
    NoC_1_24_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_1_23_io_dataIn_bits_dataType = NoC_1_24_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_1_23_io_filter_ready = pes_1_23_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_1_23_io_ifmap_ready = pes_1_23_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_1_23_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_0_clock = clock;
  assign NoC_2_0_reset = reset;
  assign NoC_2_0_io_dataPackageIn_valid = io_dataIn_valid; // @[PEArray.scala 84:35]
  assign NoC_2_0_io_dataPackageIn_bits_data = io_dataIn_bits_data; // @[PEArray.scala 85:34]
  assign NoC_2_0_io_dataPackageIn_bits_dataType = io_dataIn_bits_dataType; // @[PEArray.scala 85:34]
  assign NoC_2_0_io_dataPackageIn_bits_positon_row = io_dataIn_bits_positon_row; // @[PEArray.scala 85:34]
  assign NoC_2_0_io_dataPackageIn_bits_positon_col = io_dataIn_bits_positon_col; // @[PEArray.scala 85:34]
  assign NoC_2_0_io_dataPackageOut_ready = NoC_2_1_io_dataPackageIn_ready | NoC_2_2_io_dataPackageIn_ready |
    NoC_2_3_io_dataPackageIn_ready | NoC_2_4_io_dataPackageIn_ready | NoC_2_5_io_dataPackageIn_ready |
    NoC_2_6_io_dataPackageIn_ready | NoC_2_7_io_dataPackageIn_ready | NoC_2_8_io_dataPackageIn_ready |
    NoC_2_9_io_dataPackageIn_ready | NoC_2_10_io_dataPackageIn_ready | NoC_2_11_io_dataPackageIn_ready |
    NoC_2_12_io_dataPackageIn_ready | NoC_2_13_io_dataPackageIn_ready | NoC_2_14_io_dataPackageIn_ready |
    NoC_2_15_io_dataPackageIn_ready | NoC_2_16_io_dataPackageIn_ready | NoC_2_17_io_dataPackageIn_ready |
    NoC_2_18_io_dataPackageIn_ready | NoC_2_19_io_dataPackageIn_ready | NoC_2_20_io_dataPackageIn_ready |
    NoC_2_21_io_dataPackageIn_ready | NoC_2_22_io_dataPackageIn_ready | NoC_2_23_io_dataPackageIn_ready |
    NoC_2_24_io_dataPackageIn_ready; // @[PEArray.scala 83:17]
  assign NoC_2_1_clock = clock;
  assign NoC_2_1_reset = reset;
  assign NoC_2_1_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_1_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_1_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_1_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_1_io_dataPackageOut_ready = dss_2_0_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_0_clock = clock;
  assign pes_2_0_reset = reset;
  assign pes_2_0_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_0_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_0_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_0_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_0_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_0_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_0_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_0_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_0_io_filter_valid = dss_2_0_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_0_io_filter_bits = dss_2_0_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_0_io_ifmap_valid = dss_2_0_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_0_io_ifmap_bits = dss_2_0_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_0_io_pSumIn_valid = pes_1_0_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_0_io_pSumIn_bits = pes_1_0_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_0_io_pSumOut_ready = io_oSumOut_0_ready; // @[PEArray.scala 53:31]
  assign dss_2_0_io_dataIn_valid = NoC_2_1_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_0_io_dataIn_bits_data = {{11{NoC_2_1_io_dataPackageOut_bits_data[4]}},NoC_2_1_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_2_0_io_dataIn_bits_dataType = NoC_2_1_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_0_io_filter_ready = pes_2_0_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_0_io_ifmap_ready = pes_2_0_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_0_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_2_clock = clock;
  assign NoC_2_2_reset = reset;
  assign NoC_2_2_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_2_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_2_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_2_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_2_io_dataPackageOut_ready = dss_2_1_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_1_clock = clock;
  assign pes_2_1_reset = reset;
  assign pes_2_1_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_1_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_1_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_1_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_1_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_1_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_1_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_1_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_1_io_filter_valid = dss_2_1_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_1_io_filter_bits = dss_2_1_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_1_io_ifmap_valid = dss_2_1_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_1_io_ifmap_bits = dss_2_1_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_1_io_pSumIn_valid = pes_1_1_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_1_io_pSumIn_bits = pes_1_1_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_1_io_pSumOut_ready = io_oSumOut_1_ready; // @[PEArray.scala 53:31]
  assign dss_2_1_io_dataIn_valid = NoC_2_2_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_1_io_dataIn_bits_data = {{11{NoC_2_2_io_dataPackageOut_bits_data[4]}},NoC_2_2_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_2_1_io_dataIn_bits_dataType = NoC_2_2_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_1_io_filter_ready = pes_2_1_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_1_io_ifmap_ready = pes_2_1_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_1_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_3_clock = clock;
  assign NoC_2_3_reset = reset;
  assign NoC_2_3_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_3_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_3_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_3_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_3_io_dataPackageOut_ready = dss_2_2_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_2_clock = clock;
  assign pes_2_2_reset = reset;
  assign pes_2_2_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_2_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_2_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_2_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_2_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_2_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_2_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_2_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_2_io_filter_valid = dss_2_2_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_2_io_filter_bits = dss_2_2_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_2_io_ifmap_valid = dss_2_2_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_2_io_ifmap_bits = dss_2_2_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_2_io_pSumIn_valid = pes_1_2_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_2_io_pSumIn_bits = pes_1_2_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_2_io_pSumOut_ready = io_oSumOut_2_ready; // @[PEArray.scala 53:31]
  assign dss_2_2_io_dataIn_valid = NoC_2_3_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_2_io_dataIn_bits_data = {{11{NoC_2_3_io_dataPackageOut_bits_data[4]}},NoC_2_3_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_2_2_io_dataIn_bits_dataType = NoC_2_3_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_2_io_filter_ready = pes_2_2_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_2_io_ifmap_ready = pes_2_2_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_2_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_4_clock = clock;
  assign NoC_2_4_reset = reset;
  assign NoC_2_4_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_4_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_4_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_4_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_4_io_dataPackageOut_ready = dss_2_3_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_3_clock = clock;
  assign pes_2_3_reset = reset;
  assign pes_2_3_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_3_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_3_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_3_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_3_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_3_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_3_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_3_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_3_io_filter_valid = dss_2_3_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_3_io_filter_bits = dss_2_3_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_3_io_ifmap_valid = dss_2_3_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_3_io_ifmap_bits = dss_2_3_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_3_io_pSumIn_valid = pes_1_3_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_3_io_pSumIn_bits = pes_1_3_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_3_io_pSumOut_ready = io_oSumOut_3_ready; // @[PEArray.scala 53:31]
  assign dss_2_3_io_dataIn_valid = NoC_2_4_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_3_io_dataIn_bits_data = {{11{NoC_2_4_io_dataPackageOut_bits_data[4]}},NoC_2_4_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_2_3_io_dataIn_bits_dataType = NoC_2_4_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_3_io_filter_ready = pes_2_3_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_3_io_ifmap_ready = pes_2_3_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_3_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_5_clock = clock;
  assign NoC_2_5_reset = reset;
  assign NoC_2_5_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_5_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_5_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_5_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_5_io_dataPackageOut_ready = dss_2_4_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_4_clock = clock;
  assign pes_2_4_reset = reset;
  assign pes_2_4_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_4_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_4_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_4_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_4_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_4_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_4_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_4_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_4_io_filter_valid = dss_2_4_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_4_io_filter_bits = dss_2_4_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_4_io_ifmap_valid = dss_2_4_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_4_io_ifmap_bits = dss_2_4_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_4_io_pSumIn_valid = pes_1_4_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_4_io_pSumIn_bits = pes_1_4_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_4_io_pSumOut_ready = io_oSumOut_4_ready; // @[PEArray.scala 53:31]
  assign dss_2_4_io_dataIn_valid = NoC_2_5_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_4_io_dataIn_bits_data = {{11{NoC_2_5_io_dataPackageOut_bits_data[4]}},NoC_2_5_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_2_4_io_dataIn_bits_dataType = NoC_2_5_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_4_io_filter_ready = pes_2_4_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_4_io_ifmap_ready = pes_2_4_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_4_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_6_clock = clock;
  assign NoC_2_6_reset = reset;
  assign NoC_2_6_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_6_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_6_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_6_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_6_io_dataPackageOut_ready = dss_2_5_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_5_clock = clock;
  assign pes_2_5_reset = reset;
  assign pes_2_5_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_5_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_5_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_5_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_5_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_5_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_5_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_5_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_5_io_filter_valid = dss_2_5_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_5_io_filter_bits = dss_2_5_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_5_io_ifmap_valid = dss_2_5_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_5_io_ifmap_bits = dss_2_5_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_5_io_pSumIn_valid = pes_1_5_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_5_io_pSumIn_bits = pes_1_5_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_5_io_pSumOut_ready = io_oSumOut_5_ready; // @[PEArray.scala 53:31]
  assign dss_2_5_io_dataIn_valid = NoC_2_6_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_5_io_dataIn_bits_data = {{11{NoC_2_6_io_dataPackageOut_bits_data[4]}},NoC_2_6_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_2_5_io_dataIn_bits_dataType = NoC_2_6_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_5_io_filter_ready = pes_2_5_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_5_io_ifmap_ready = pes_2_5_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_5_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_7_clock = clock;
  assign NoC_2_7_reset = reset;
  assign NoC_2_7_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_7_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_7_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_7_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_7_io_dataPackageOut_ready = dss_2_6_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_6_clock = clock;
  assign pes_2_6_reset = reset;
  assign pes_2_6_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_6_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_6_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_6_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_6_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_6_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_6_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_6_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_6_io_filter_valid = dss_2_6_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_6_io_filter_bits = dss_2_6_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_6_io_ifmap_valid = dss_2_6_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_6_io_ifmap_bits = dss_2_6_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_6_io_pSumIn_valid = pes_1_6_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_6_io_pSumIn_bits = pes_1_6_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_6_io_pSumOut_ready = io_oSumOut_6_ready; // @[PEArray.scala 53:31]
  assign dss_2_6_io_dataIn_valid = NoC_2_7_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_6_io_dataIn_bits_data = {{11{NoC_2_7_io_dataPackageOut_bits_data[4]}},NoC_2_7_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_2_6_io_dataIn_bits_dataType = NoC_2_7_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_6_io_filter_ready = pes_2_6_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_6_io_ifmap_ready = pes_2_6_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_6_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_8_clock = clock;
  assign NoC_2_8_reset = reset;
  assign NoC_2_8_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_8_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_8_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_8_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_8_io_dataPackageOut_ready = dss_2_7_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_7_clock = clock;
  assign pes_2_7_reset = reset;
  assign pes_2_7_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_7_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_7_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_7_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_7_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_7_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_7_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_7_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_7_io_filter_valid = dss_2_7_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_7_io_filter_bits = dss_2_7_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_7_io_ifmap_valid = dss_2_7_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_7_io_ifmap_bits = dss_2_7_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_7_io_pSumIn_valid = pes_1_7_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_7_io_pSumIn_bits = pes_1_7_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_7_io_pSumOut_ready = io_oSumOut_7_ready; // @[PEArray.scala 53:31]
  assign dss_2_7_io_dataIn_valid = NoC_2_8_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_7_io_dataIn_bits_data = {{11{NoC_2_8_io_dataPackageOut_bits_data[4]}},NoC_2_8_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_2_7_io_dataIn_bits_dataType = NoC_2_8_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_7_io_filter_ready = pes_2_7_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_7_io_ifmap_ready = pes_2_7_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_7_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_9_clock = clock;
  assign NoC_2_9_reset = reset;
  assign NoC_2_9_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_9_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_9_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_9_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_9_io_dataPackageOut_ready = dss_2_8_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_8_clock = clock;
  assign pes_2_8_reset = reset;
  assign pes_2_8_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_8_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_8_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_8_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_8_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_8_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_8_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_8_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_8_io_filter_valid = dss_2_8_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_8_io_filter_bits = dss_2_8_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_8_io_ifmap_valid = dss_2_8_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_8_io_ifmap_bits = dss_2_8_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_8_io_pSumIn_valid = pes_1_8_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_8_io_pSumIn_bits = pes_1_8_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_8_io_pSumOut_ready = io_oSumOut_8_ready; // @[PEArray.scala 53:31]
  assign dss_2_8_io_dataIn_valid = NoC_2_9_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_8_io_dataIn_bits_data = {{11{NoC_2_9_io_dataPackageOut_bits_data[4]}},NoC_2_9_io_dataPackageOut_bits_data
    }; // @[PEArray.scala 38:22]
  assign dss_2_8_io_dataIn_bits_dataType = NoC_2_9_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_8_io_filter_ready = pes_2_8_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_8_io_ifmap_ready = pes_2_8_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_8_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_10_clock = clock;
  assign NoC_2_10_reset = reset;
  assign NoC_2_10_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_10_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_10_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_10_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_10_io_dataPackageOut_ready = dss_2_9_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_9_clock = clock;
  assign pes_2_9_reset = reset;
  assign pes_2_9_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_9_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_9_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_9_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_9_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_9_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_9_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_9_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_9_io_filter_valid = dss_2_9_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_9_io_filter_bits = dss_2_9_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_9_io_ifmap_valid = dss_2_9_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_9_io_ifmap_bits = dss_2_9_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_9_io_pSumIn_valid = pes_1_9_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_9_io_pSumIn_bits = pes_1_9_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_9_io_pSumOut_ready = io_oSumOut_9_ready; // @[PEArray.scala 53:31]
  assign dss_2_9_io_dataIn_valid = NoC_2_10_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_9_io_dataIn_bits_data = {{11{NoC_2_10_io_dataPackageOut_bits_data[4]}},
    NoC_2_10_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_9_io_dataIn_bits_dataType = NoC_2_10_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_9_io_filter_ready = pes_2_9_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_9_io_ifmap_ready = pes_2_9_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_9_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_11_clock = clock;
  assign NoC_2_11_reset = reset;
  assign NoC_2_11_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_11_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_11_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_11_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_11_io_dataPackageOut_ready = dss_2_10_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_10_clock = clock;
  assign pes_2_10_reset = reset;
  assign pes_2_10_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_10_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_10_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_10_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_10_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_10_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_10_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_10_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_10_io_filter_valid = dss_2_10_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_10_io_filter_bits = dss_2_10_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_10_io_ifmap_valid = dss_2_10_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_10_io_ifmap_bits = dss_2_10_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_10_io_pSumIn_valid = pes_1_10_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_10_io_pSumIn_bits = pes_1_10_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_10_io_pSumOut_ready = io_oSumOut_10_ready; // @[PEArray.scala 53:31]
  assign dss_2_10_io_dataIn_valid = NoC_2_11_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_10_io_dataIn_bits_data = {{11{NoC_2_11_io_dataPackageOut_bits_data[4]}},
    NoC_2_11_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_10_io_dataIn_bits_dataType = NoC_2_11_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_10_io_filter_ready = pes_2_10_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_10_io_ifmap_ready = pes_2_10_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_10_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_12_clock = clock;
  assign NoC_2_12_reset = reset;
  assign NoC_2_12_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_12_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_12_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_12_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_12_io_dataPackageOut_ready = dss_2_11_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_11_clock = clock;
  assign pes_2_11_reset = reset;
  assign pes_2_11_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_11_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_11_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_11_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_11_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_11_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_11_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_11_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_11_io_filter_valid = dss_2_11_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_11_io_filter_bits = dss_2_11_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_11_io_ifmap_valid = dss_2_11_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_11_io_ifmap_bits = dss_2_11_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_11_io_pSumIn_valid = pes_1_11_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_11_io_pSumIn_bits = pes_1_11_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_11_io_pSumOut_ready = io_oSumOut_11_ready; // @[PEArray.scala 53:31]
  assign dss_2_11_io_dataIn_valid = NoC_2_12_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_11_io_dataIn_bits_data = {{11{NoC_2_12_io_dataPackageOut_bits_data[4]}},
    NoC_2_12_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_11_io_dataIn_bits_dataType = NoC_2_12_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_11_io_filter_ready = pes_2_11_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_11_io_ifmap_ready = pes_2_11_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_11_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_13_clock = clock;
  assign NoC_2_13_reset = reset;
  assign NoC_2_13_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_13_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_13_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_13_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_13_io_dataPackageOut_ready = dss_2_12_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_12_clock = clock;
  assign pes_2_12_reset = reset;
  assign pes_2_12_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_12_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_12_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_12_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_12_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_12_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_12_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_12_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_12_io_filter_valid = dss_2_12_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_12_io_filter_bits = dss_2_12_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_12_io_ifmap_valid = dss_2_12_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_12_io_ifmap_bits = dss_2_12_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_12_io_pSumIn_valid = pes_1_12_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_12_io_pSumIn_bits = pes_1_12_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_12_io_pSumOut_ready = io_oSumOut_12_ready; // @[PEArray.scala 53:31]
  assign dss_2_12_io_dataIn_valid = NoC_2_13_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_12_io_dataIn_bits_data = {{11{NoC_2_13_io_dataPackageOut_bits_data[4]}},
    NoC_2_13_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_12_io_dataIn_bits_dataType = NoC_2_13_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_12_io_filter_ready = pes_2_12_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_12_io_ifmap_ready = pes_2_12_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_12_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_14_clock = clock;
  assign NoC_2_14_reset = reset;
  assign NoC_2_14_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_14_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_14_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_14_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_14_io_dataPackageOut_ready = dss_2_13_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_13_clock = clock;
  assign pes_2_13_reset = reset;
  assign pes_2_13_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_13_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_13_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_13_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_13_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_13_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_13_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_13_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_13_io_filter_valid = dss_2_13_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_13_io_filter_bits = dss_2_13_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_13_io_ifmap_valid = dss_2_13_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_13_io_ifmap_bits = dss_2_13_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_13_io_pSumIn_valid = pes_1_13_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_13_io_pSumIn_bits = pes_1_13_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_13_io_pSumOut_ready = io_oSumOut_13_ready; // @[PEArray.scala 53:31]
  assign dss_2_13_io_dataIn_valid = NoC_2_14_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_13_io_dataIn_bits_data = {{11{NoC_2_14_io_dataPackageOut_bits_data[4]}},
    NoC_2_14_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_13_io_dataIn_bits_dataType = NoC_2_14_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_13_io_filter_ready = pes_2_13_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_13_io_ifmap_ready = pes_2_13_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_13_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_15_clock = clock;
  assign NoC_2_15_reset = reset;
  assign NoC_2_15_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_15_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_15_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_15_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_15_io_dataPackageOut_ready = dss_2_14_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_14_clock = clock;
  assign pes_2_14_reset = reset;
  assign pes_2_14_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_14_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_14_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_14_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_14_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_14_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_14_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_14_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_14_io_filter_valid = dss_2_14_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_14_io_filter_bits = dss_2_14_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_14_io_ifmap_valid = dss_2_14_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_14_io_ifmap_bits = dss_2_14_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_14_io_pSumIn_valid = pes_1_14_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_14_io_pSumIn_bits = pes_1_14_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_14_io_pSumOut_ready = io_oSumOut_14_ready; // @[PEArray.scala 53:31]
  assign dss_2_14_io_dataIn_valid = NoC_2_15_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_14_io_dataIn_bits_data = {{11{NoC_2_15_io_dataPackageOut_bits_data[4]}},
    NoC_2_15_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_14_io_dataIn_bits_dataType = NoC_2_15_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_14_io_filter_ready = pes_2_14_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_14_io_ifmap_ready = pes_2_14_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_14_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_16_clock = clock;
  assign NoC_2_16_reset = reset;
  assign NoC_2_16_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_16_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_16_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_16_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_16_io_dataPackageOut_ready = dss_2_15_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_15_clock = clock;
  assign pes_2_15_reset = reset;
  assign pes_2_15_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_15_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_15_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_15_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_15_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_15_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_15_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_15_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_15_io_filter_valid = dss_2_15_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_15_io_filter_bits = dss_2_15_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_15_io_ifmap_valid = dss_2_15_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_15_io_ifmap_bits = dss_2_15_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_15_io_pSumIn_valid = pes_1_15_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_15_io_pSumIn_bits = pes_1_15_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_15_io_pSumOut_ready = io_oSumOut_15_ready; // @[PEArray.scala 53:31]
  assign dss_2_15_io_dataIn_valid = NoC_2_16_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_15_io_dataIn_bits_data = {{11{NoC_2_16_io_dataPackageOut_bits_data[4]}},
    NoC_2_16_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_15_io_dataIn_bits_dataType = NoC_2_16_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_15_io_filter_ready = pes_2_15_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_15_io_ifmap_ready = pes_2_15_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_15_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_17_clock = clock;
  assign NoC_2_17_reset = reset;
  assign NoC_2_17_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_17_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_17_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_17_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_17_io_dataPackageOut_ready = dss_2_16_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_16_clock = clock;
  assign pes_2_16_reset = reset;
  assign pes_2_16_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_16_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_16_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_16_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_16_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_16_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_16_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_16_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_16_io_filter_valid = dss_2_16_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_16_io_filter_bits = dss_2_16_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_16_io_ifmap_valid = dss_2_16_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_16_io_ifmap_bits = dss_2_16_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_16_io_pSumIn_valid = pes_1_16_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_16_io_pSumIn_bits = pes_1_16_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_16_io_pSumOut_ready = io_oSumOut_16_ready; // @[PEArray.scala 53:31]
  assign dss_2_16_io_dataIn_valid = NoC_2_17_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_16_io_dataIn_bits_data = {{11{NoC_2_17_io_dataPackageOut_bits_data[4]}},
    NoC_2_17_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_16_io_dataIn_bits_dataType = NoC_2_17_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_16_io_filter_ready = pes_2_16_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_16_io_ifmap_ready = pes_2_16_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_16_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_18_clock = clock;
  assign NoC_2_18_reset = reset;
  assign NoC_2_18_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_18_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_18_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_18_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_18_io_dataPackageOut_ready = dss_2_17_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_17_clock = clock;
  assign pes_2_17_reset = reset;
  assign pes_2_17_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_17_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_17_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_17_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_17_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_17_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_17_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_17_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_17_io_filter_valid = dss_2_17_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_17_io_filter_bits = dss_2_17_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_17_io_ifmap_valid = dss_2_17_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_17_io_ifmap_bits = dss_2_17_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_17_io_pSumIn_valid = pes_1_17_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_17_io_pSumIn_bits = pes_1_17_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_17_io_pSumOut_ready = io_oSumOut_17_ready; // @[PEArray.scala 53:31]
  assign dss_2_17_io_dataIn_valid = NoC_2_18_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_17_io_dataIn_bits_data = {{11{NoC_2_18_io_dataPackageOut_bits_data[4]}},
    NoC_2_18_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_17_io_dataIn_bits_dataType = NoC_2_18_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_17_io_filter_ready = pes_2_17_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_17_io_ifmap_ready = pes_2_17_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_17_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_19_clock = clock;
  assign NoC_2_19_reset = reset;
  assign NoC_2_19_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_19_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_19_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_19_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_19_io_dataPackageOut_ready = dss_2_18_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_18_clock = clock;
  assign pes_2_18_reset = reset;
  assign pes_2_18_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_18_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_18_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_18_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_18_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_18_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_18_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_18_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_18_io_filter_valid = dss_2_18_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_18_io_filter_bits = dss_2_18_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_18_io_ifmap_valid = dss_2_18_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_18_io_ifmap_bits = dss_2_18_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_18_io_pSumIn_valid = pes_1_18_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_18_io_pSumIn_bits = pes_1_18_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_18_io_pSumOut_ready = io_oSumOut_18_ready; // @[PEArray.scala 53:31]
  assign dss_2_18_io_dataIn_valid = NoC_2_19_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_18_io_dataIn_bits_data = {{11{NoC_2_19_io_dataPackageOut_bits_data[4]}},
    NoC_2_19_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_18_io_dataIn_bits_dataType = NoC_2_19_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_18_io_filter_ready = pes_2_18_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_18_io_ifmap_ready = pes_2_18_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_18_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_20_clock = clock;
  assign NoC_2_20_reset = reset;
  assign NoC_2_20_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_20_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_20_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_20_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_20_io_dataPackageOut_ready = dss_2_19_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_19_clock = clock;
  assign pes_2_19_reset = reset;
  assign pes_2_19_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_19_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_19_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_19_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_19_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_19_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_19_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_19_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_19_io_filter_valid = dss_2_19_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_19_io_filter_bits = dss_2_19_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_19_io_ifmap_valid = dss_2_19_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_19_io_ifmap_bits = dss_2_19_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_19_io_pSumIn_valid = pes_1_19_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_19_io_pSumIn_bits = pes_1_19_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_19_io_pSumOut_ready = io_oSumOut_19_ready; // @[PEArray.scala 53:31]
  assign dss_2_19_io_dataIn_valid = NoC_2_20_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_19_io_dataIn_bits_data = {{11{NoC_2_20_io_dataPackageOut_bits_data[4]}},
    NoC_2_20_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_19_io_dataIn_bits_dataType = NoC_2_20_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_19_io_filter_ready = pes_2_19_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_19_io_ifmap_ready = pes_2_19_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_19_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_21_clock = clock;
  assign NoC_2_21_reset = reset;
  assign NoC_2_21_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_21_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_21_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_21_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_21_io_dataPackageOut_ready = dss_2_20_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_20_clock = clock;
  assign pes_2_20_reset = reset;
  assign pes_2_20_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_20_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_20_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_20_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_20_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_20_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_20_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_20_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_20_io_filter_valid = dss_2_20_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_20_io_filter_bits = dss_2_20_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_20_io_ifmap_valid = dss_2_20_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_20_io_ifmap_bits = dss_2_20_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_20_io_pSumIn_valid = pes_1_20_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_20_io_pSumIn_bits = pes_1_20_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_20_io_pSumOut_ready = io_oSumOut_20_ready; // @[PEArray.scala 53:31]
  assign dss_2_20_io_dataIn_valid = NoC_2_21_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_20_io_dataIn_bits_data = {{11{NoC_2_21_io_dataPackageOut_bits_data[4]}},
    NoC_2_21_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_20_io_dataIn_bits_dataType = NoC_2_21_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_20_io_filter_ready = pes_2_20_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_20_io_ifmap_ready = pes_2_20_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_20_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_22_clock = clock;
  assign NoC_2_22_reset = reset;
  assign NoC_2_22_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_22_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_22_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_22_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_22_io_dataPackageOut_ready = dss_2_21_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_21_clock = clock;
  assign pes_2_21_reset = reset;
  assign pes_2_21_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_21_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_21_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_21_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_21_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_21_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_21_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_21_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_21_io_filter_valid = dss_2_21_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_21_io_filter_bits = dss_2_21_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_21_io_ifmap_valid = dss_2_21_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_21_io_ifmap_bits = dss_2_21_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_21_io_pSumIn_valid = pes_1_21_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_21_io_pSumIn_bits = pes_1_21_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_21_io_pSumOut_ready = io_oSumOut_21_ready; // @[PEArray.scala 53:31]
  assign dss_2_21_io_dataIn_valid = NoC_2_22_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_21_io_dataIn_bits_data = {{11{NoC_2_22_io_dataPackageOut_bits_data[4]}},
    NoC_2_22_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_21_io_dataIn_bits_dataType = NoC_2_22_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_21_io_filter_ready = pes_2_21_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_21_io_ifmap_ready = pes_2_21_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_21_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_23_clock = clock;
  assign NoC_2_23_reset = reset;
  assign NoC_2_23_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_23_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_23_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_23_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_23_io_dataPackageOut_ready = dss_2_22_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_22_clock = clock;
  assign pes_2_22_reset = reset;
  assign pes_2_22_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_22_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_22_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_22_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_22_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_22_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_22_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_22_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_22_io_filter_valid = dss_2_22_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_22_io_filter_bits = dss_2_22_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_22_io_ifmap_valid = dss_2_22_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_22_io_ifmap_bits = dss_2_22_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_22_io_pSumIn_valid = pes_1_22_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_22_io_pSumIn_bits = pes_1_22_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_22_io_pSumOut_ready = io_oSumOut_22_ready; // @[PEArray.scala 53:31]
  assign dss_2_22_io_dataIn_valid = NoC_2_23_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_22_io_dataIn_bits_data = {{11{NoC_2_23_io_dataPackageOut_bits_data[4]}},
    NoC_2_23_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_22_io_dataIn_bits_dataType = NoC_2_23_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_22_io_filter_ready = pes_2_22_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_22_io_ifmap_ready = pes_2_22_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_22_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  assign NoC_2_24_clock = clock;
  assign NoC_2_24_reset = reset;
  assign NoC_2_24_io_dataPackageIn_valid = NoC_2_0_io_dataPackageOut_valid; // @[PEArray.scala 74:40]
  assign NoC_2_24_io_dataPackageIn_bits_data = NoC_2_0_io_dataPackageOut_bits_data; // @[PEArray.scala 75:39]
  assign NoC_2_24_io_dataPackageIn_bits_dataType = NoC_2_0_io_dataPackageOut_bits_dataType; // @[PEArray.scala 75:39]
  assign NoC_2_24_io_dataPackageIn_bits_positon_col = NoC_2_0_io_dataPackageOut_bits_positon_col; // @[PEArray.scala 75:39]
  assign NoC_2_24_io_dataPackageOut_ready = dss_2_23_io_dataIn_ready; // @[PEArray.scala 38:22]
  assign pes_2_23_clock = clock;
  assign pes_2_23_reset = reset;
  assign pes_2_23_io_stateSW = io_stateSW; // @[PEArray.scala 44:23]
  assign pes_2_23_io_peconfig_valid = io_peconfig_valid; // @[PEArray.scala 43:30]
  assign pes_2_23_io_peconfig_bits_ichannelNum = io_peconfig_bits_ichannelNum; // @[PEArray.scala 42:29]
  assign pes_2_23_io_peconfig_bits_ochannelNum = io_peconfig_bits_ochannelNum; // @[PEArray.scala 42:29]
  assign pes_2_23_io_peconfig_bits_ofmapW = io_peconfig_bits_ofmapW; // @[PEArray.scala 42:29]
  assign pes_2_23_io_peconfig_bits_stepW = io_peconfig_bits_stepW; // @[PEArray.scala 42:29]
  assign pes_2_23_io_peconfig_bits_filterLen = io_peconfig_bits_filterLen; // @[PEArray.scala 42:29]
  assign pes_2_23_io_peconfig_bits_ifmapLen = io_peconfig_bits_ifmapLen; // @[PEArray.scala 42:29]
  assign pes_2_23_io_filter_valid = dss_2_23_io_filter_valid; // @[PEArray.scala 39:22]
  assign pes_2_23_io_filter_bits = dss_2_23_io_filter_bits[4:0]; // @[PEArray.scala 39:22]
  assign pes_2_23_io_ifmap_valid = dss_2_23_io_ifmap_valid; // @[PEArray.scala 40:21]
  assign pes_2_23_io_ifmap_bits = dss_2_23_io_ifmap_bits[4:0]; // @[PEArray.scala 40:21]
  assign pes_2_23_io_pSumIn_valid = pes_1_23_io_pSumOut_valid; // @[PEArray.scala 93:27]
  assign pes_2_23_io_pSumIn_bits = pes_1_23_io_pSumOut_bits; // @[PEArray.scala 93:27]
  assign pes_2_23_io_pSumOut_ready = io_oSumOut_23_ready; // @[PEArray.scala 53:31]
  assign dss_2_23_io_dataIn_valid = NoC_2_24_io_dataPackageOut_valid; // @[PEArray.scala 38:22]
  assign dss_2_23_io_dataIn_bits_data = {{11{NoC_2_24_io_dataPackageOut_bits_data[4]}},
    NoC_2_24_io_dataPackageOut_bits_data}; // @[PEArray.scala 38:22]
  assign dss_2_23_io_dataIn_bits_dataType = NoC_2_24_io_dataPackageOut_bits_dataType; // @[PEArray.scala 38:22]
  assign dss_2_23_io_filter_ready = pes_2_23_io_filter_ready; // @[PEArray.scala 39:22]
  assign dss_2_23_io_ifmap_ready = pes_2_23_io_ifmap_ready; // @[PEArray.scala 40:21]
  assign dss_2_23_io_pSum_ready = 1'h0; // @[PEArray.scala 48:28]
  always @(posedge clock) begin
    if (reset) begin // @[PEArray.scala 17:24]
      doneReg <= 1'h0; // @[PEArray.scala 17:24]
    end else begin
      doneReg <= _T_182 | pes_2_16_io_stateOut == 4'h6 | pes_2_17_io_stateOut == 4'h6 | pes_2_18_io_stateOut == 4'h6 |
        pes_2_19_io_stateOut == 4'h6 | pes_2_20_io_stateOut == 4'h6 | pes_2_21_io_stateOut == 4'h6 |
        pes_2_22_io_stateOut == 4'h6 | pes_2_23_io_stateOut == 4'h6; // @[PEArray.scala 103:11]
    end
    if (_T) begin // @[PEArray.scala 21:28]
      configReg_relu <= io_peconfig_bits_relu; // @[PEArray.scala 22:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  doneReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  configReg_relu = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
